*-- interposer PDN spice model 'interposer' for AC analysis
*-- Total unit cell #: 121 (11x11)

.param cellno=121
.param r_int_cell='1e-3'
.param l_int_cell='1e-10'
.param c_int_cell='1e-11'

xdint_0_0 ndint_x_0_0 ndint_x_909_0 ndint_y_0_0 ndint_y_0_909 ndint_xy_0_0 int_unitcell rval='r_int_cell' lval='l_int_cell' cval='c_int_cell'
xdint_0_1 ndint_x_909_0 ndint_x_1818_0 ndint_y_909_0 ndint_y_909_909 ndint_xy_909_0 int_unitcell rval='r_int_cell' lval='l_int_cell' cval='c_int_cell'
xdint_0_2 ndint_x_1818_0 ndint_x_2727_0 ndint_y_1818_0 ndint_y_1818_909 ndint_xy_1818_0 int_unitcell rval='r_int_cell' lval='l_int_cell' cval='c_int_cell'
xdint_0_3 ndint_x_2727_0 ndint_x_3636_0 ndint_y_2727_0 ndint_y_2727_909 ndint_xy_2727_0 int_unitcell rval='r_int_cell' lval='l_int_cell' cval='c_int_cell'
xdint_0_4 ndint_x_3636_0 ndint_x_4545_0 ndint_y_3636_0 ndint_y_3636_909 ndint_xy_3636_0 int_unitcell rval='r_int_cell' lval='l_int_cell' cval='c_int_cell'
xdint_0_5 ndint_x_4545_0 ndint_x_5454_0 ndint_y_4545_0 ndint_y_4545_909 ndint_xy_4545_0 int_unitcell rval='r_int_cell' lval='l_int_cell' cval='c_int_cell'
xdint_0_6 ndint_x_5454_0 ndint_x_6363_0 ndint_y_5454_0 ndint_y_5454_909 ndint_xy_5454_0 int_unitcell rval='r_int_cell' lval='l_int_cell' cval='c_int_cell'
xdint_0_7 ndint_x_6363_0 ndint_x_7272_0 ndint_y_6363_0 ndint_y_6363_909 ndint_xy_6363_0 int_unitcell rval='r_int_cell' lval='l_int_cell' cval='c_int_cell'
xdint_0_8 ndint_x_7272_0 ndint_x_8181_0 ndint_y_7272_0 ndint_y_7272_909 ndint_xy_7272_0 int_unitcell rval='r_int_cell' lval='l_int_cell' cval='c_int_cell'
xdint_0_9 ndint_x_8181_0 ndint_x_9090_0 ndint_y_8181_0 ndint_y_8181_909 ndint_xy_8181_0 int_unitcell rval='r_int_cell' lval='l_int_cell' cval='c_int_cell'
xdint_0_10 ndint_x_9090_0 ndint_x_9999_0 ndint_y_9090_0 ndint_y_9090_909 ndint_xy_9090_0 int_unitcell rval='r_int_cell' lval='l_int_cell' cval='c_int_cell'
xdint_1_0 ndint_x_0_909 ndint_x_909_909 ndint_y_0_909 ndint_y_0_1818 ndint_xy_0_909 int_unitcell rval='r_int_cell' lval='l_int_cell' cval='c_int_cell'
xdint_1_1 ndint_x_909_909 ndint_x_1818_909 ndint_y_909_909 ndint_y_909_1818 ndint_xy_909_909 int_unitcell rval='r_int_cell' lval='l_int_cell' cval='c_int_cell'
xdint_1_2 ndint_x_1818_909 ndint_x_2727_909 ndint_y_1818_909 ndint_y_1818_1818 ndint_xy_1818_909 int_unitcell rval='r_int_cell' lval='l_int_cell' cval='c_int_cell'
xdint_1_3 ndint_x_2727_909 ndint_x_3636_909 ndint_y_2727_909 ndint_y_2727_1818 ndint_xy_2727_909 int_unitcell rval='r_int_cell' lval='l_int_cell' cval='c_int_cell'
xdint_1_4 ndint_x_3636_909 ndint_x_4545_909 ndint_y_3636_909 ndint_y_3636_1818 ndint_xy_3636_909 int_unitcell rval='r_int_cell' lval='l_int_cell' cval='c_int_cell'
xdint_1_5 ndint_x_4545_909 ndint_x_5454_909 ndint_y_4545_909 ndint_y_4545_1818 ndint_xy_4545_909 int_unitcell rval='r_int_cell' lval='l_int_cell' cval='c_int_cell'
xdint_1_6 ndint_x_5454_909 ndint_x_6363_909 ndint_y_5454_909 ndint_y_5454_1818 ndint_xy_5454_909 int_unitcell rval='r_int_cell' lval='l_int_cell' cval='c_int_cell'
xdint_1_7 ndint_x_6363_909 ndint_x_7272_909 ndint_y_6363_909 ndint_y_6363_1818 ndint_xy_6363_909 int_unitcell rval='r_int_cell' lval='l_int_cell' cval='c_int_cell'
xdint_1_8 ndint_x_7272_909 ndint_x_8181_909 ndint_y_7272_909 ndint_y_7272_1818 ndint_xy_7272_909 int_unitcell rval='r_int_cell' lval='l_int_cell' cval='c_int_cell'
xdint_1_9 ndint_x_8181_909 ndint_x_9090_909 ndint_y_8181_909 ndint_y_8181_1818 ndint_xy_8181_909 int_unitcell rval='r_int_cell' lval='l_int_cell' cval='c_int_cell'
xdint_1_10 ndint_x_9090_909 ndint_x_9999_909 ndint_y_9090_909 ndint_y_9090_1818 ndint_xy_9090_909 int_unitcell rval='r_int_cell' lval='l_int_cell' cval='c_int_cell'
xdint_2_0 ndint_x_0_1818 ndint_x_909_1818 ndint_y_0_1818 ndint_y_0_2727 ndint_xy_0_1818 int_unitcell rval='r_int_cell' lval='l_int_cell' cval='c_int_cell'
xdint_2_1 ndint_x_909_1818 ndint_x_1818_1818 ndint_y_909_1818 ndint_y_909_2727 ndint_xy_909_1818 int_unitcell rval='r_int_cell' lval='l_int_cell' cval='c_int_cell'
xdint_2_2 ndint_x_1818_1818 ndint_x_2727_1818 ndint_y_1818_1818 ndint_y_1818_2727 ndint_xy_1818_1818 int_unitcell rval='r_int_cell' lval='l_int_cell' cval='c_int_cell'
xdint_2_3 ndint_x_2727_1818 ndint_x_3636_1818 ndint_y_2727_1818 ndint_y_2727_2727 ndint_xy_2727_1818 int_unitcell rval='r_int_cell' lval='l_int_cell' cval='c_int_cell'
xdint_2_4 ndint_x_3636_1818 ndint_x_4545_1818 ndint_y_3636_1818 ndint_y_3636_2727 ndint_xy_3636_1818 int_unitcell rval='r_int_cell' lval='l_int_cell' cval='c_int_cell'
xdint_2_5 ndint_x_4545_1818 ndint_x_5454_1818 ndint_y_4545_1818 ndint_y_4545_2727 ndint_xy_4545_1818 int_unitcell rval='r_int_cell' lval='l_int_cell' cval='c_int_cell'
xdint_2_6 ndint_x_5454_1818 ndint_x_6363_1818 ndint_y_5454_1818 ndint_y_5454_2727 ndint_xy_5454_1818 int_unitcell rval='r_int_cell' lval='l_int_cell' cval='c_int_cell'
xdint_2_7 ndint_x_6363_1818 ndint_x_7272_1818 ndint_y_6363_1818 ndint_y_6363_2727 ndint_xy_6363_1818 int_unitcell rval='r_int_cell' lval='l_int_cell' cval='c_int_cell'
xdint_2_8 ndint_x_7272_1818 ndint_x_8181_1818 ndint_y_7272_1818 ndint_y_7272_2727 ndint_xy_7272_1818 int_unitcell rval='r_int_cell' lval='l_int_cell' cval='c_int_cell'
xdint_2_9 ndint_x_8181_1818 ndint_x_9090_1818 ndint_y_8181_1818 ndint_y_8181_2727 ndint_xy_8181_1818 int_unitcell rval='r_int_cell' lval='l_int_cell' cval='c_int_cell'
xdint_2_10 ndint_x_9090_1818 ndint_x_9999_1818 ndint_y_9090_1818 ndint_y_9090_2727 ndint_xy_9090_1818 int_unitcell rval='r_int_cell' lval='l_int_cell' cval='c_int_cell'
xdint_3_0 ndint_x_0_2727 ndint_x_909_2727 ndint_y_0_2727 ndint_y_0_3636 ndint_xy_0_2727 int_unitcell rval='r_int_cell' lval='l_int_cell' cval='c_int_cell'
xdint_3_1 ndint_x_909_2727 ndint_x_1818_2727 ndint_y_909_2727 ndint_y_909_3636 ndint_xy_909_2727 int_unitcell rval='r_int_cell' lval='l_int_cell' cval='c_int_cell'
xdint_3_2 ndint_x_1818_2727 ndint_x_2727_2727 ndint_y_1818_2727 ndint_y_1818_3636 ndint_xy_1818_2727 int_unitcell rval='r_int_cell' lval='l_int_cell' cval='c_int_cell'
xdint_3_3 ndint_x_2727_2727 ndint_x_3636_2727 ndint_y_2727_2727 ndint_y_2727_3636 ndint_xy_2727_2727 int_unitcell rval='r_int_cell' lval='l_int_cell' cval='c_int_cell'
xdint_3_4 ndint_x_3636_2727 ndint_x_4545_2727 ndint_y_3636_2727 ndint_y_3636_3636 ndint_xy_3636_2727 int_unitcell rval='r_int_cell' lval='l_int_cell' cval='c_int_cell'
xdint_3_5 ndint_x_4545_2727 ndint_x_5454_2727 ndint_y_4545_2727 ndint_y_4545_3636 ndint_xy_4545_2727 int_unitcell rval='r_int_cell' lval='l_int_cell' cval='c_int_cell'
xdint_3_6 ndint_x_5454_2727 ndint_x_6363_2727 ndint_y_5454_2727 ndint_y_5454_3636 ndint_xy_5454_2727 int_unitcell rval='r_int_cell' lval='l_int_cell' cval='c_int_cell'
xdint_3_7 ndint_x_6363_2727 ndint_x_7272_2727 ndint_y_6363_2727 ndint_y_6363_3636 ndint_xy_6363_2727 int_unitcell rval='r_int_cell' lval='l_int_cell' cval='c_int_cell'
xdint_3_8 ndint_x_7272_2727 ndint_x_8181_2727 ndint_y_7272_2727 ndint_y_7272_3636 ndint_xy_7272_2727 int_unitcell rval='r_int_cell' lval='l_int_cell' cval='c_int_cell'
xdint_3_9 ndint_x_8181_2727 ndint_x_9090_2727 ndint_y_8181_2727 ndint_y_8181_3636 ndint_xy_8181_2727 int_unitcell rval='r_int_cell' lval='l_int_cell' cval='c_int_cell'
xdint_3_10 ndint_x_9090_2727 ndint_x_9999_2727 ndint_y_9090_2727 ndint_y_9090_3636 ndint_xy_9090_2727 int_unitcell rval='r_int_cell' lval='l_int_cell' cval='c_int_cell'
xdint_4_0 ndint_x_0_3636 ndint_x_909_3636 ndint_y_0_3636 ndint_y_0_4545 ndint_xy_0_3636 int_unitcell rval='r_int_cell' lval='l_int_cell' cval='c_int_cell'
xdint_4_1 ndint_x_909_3636 ndint_x_1818_3636 ndint_y_909_3636 ndint_y_909_4545 ndint_xy_909_3636 int_unitcell rval='r_int_cell' lval='l_int_cell' cval='c_int_cell'
xdint_4_2 ndint_x_1818_3636 ndint_x_2727_3636 ndint_y_1818_3636 ndint_y_1818_4545 ndint_xy_1818_3636 int_unitcell rval='r_int_cell' lval='l_int_cell' cval='c_int_cell'
xdint_4_3 ndint_x_2727_3636 ndint_x_3636_3636 ndint_y_2727_3636 ndint_y_2727_4545 ndint_xy_2727_3636 int_unitcell rval='r_int_cell' lval='l_int_cell' cval='c_int_cell'
xdint_4_4 ndint_x_3636_3636 ndint_x_4545_3636 ndint_y_3636_3636 ndint_y_3636_4545 ndint_xy_3636_3636 int_unitcell rval='r_int_cell' lval='l_int_cell' cval='c_int_cell'
xdint_4_5 ndint_x_4545_3636 ndint_x_5454_3636 ndint_y_4545_3636 ndint_y_4545_4545 ndint_xy_4545_3636 int_unitcell rval='r_int_cell' lval='l_int_cell' cval='c_int_cell'
xdint_4_6 ndint_x_5454_3636 ndint_x_6363_3636 ndint_y_5454_3636 ndint_y_5454_4545 ndint_xy_5454_3636 int_unitcell rval='r_int_cell' lval='l_int_cell' cval='c_int_cell'
xdint_4_7 ndint_x_6363_3636 ndint_x_7272_3636 ndint_y_6363_3636 ndint_y_6363_4545 ndint_xy_6363_3636 int_unitcell rval='r_int_cell' lval='l_int_cell' cval='c_int_cell'
xdint_4_8 ndint_x_7272_3636 ndint_x_8181_3636 ndint_y_7272_3636 ndint_y_7272_4545 ndint_xy_7272_3636 int_unitcell rval='r_int_cell' lval='l_int_cell' cval='c_int_cell'
xdint_4_9 ndint_x_8181_3636 ndint_x_9090_3636 ndint_y_8181_3636 ndint_y_8181_4545 ndint_xy_8181_3636 int_unitcell rval='r_int_cell' lval='l_int_cell' cval='c_int_cell'
xdint_4_10 ndint_x_9090_3636 ndint_x_9999_3636 ndint_y_9090_3636 ndint_y_9090_4545 ndint_xy_9090_3636 int_unitcell rval='r_int_cell' lval='l_int_cell' cval='c_int_cell'
xdint_5_0 ndint_x_0_4545 ndint_x_909_4545 ndint_y_0_4545 ndint_y_0_5454 ndint_xy_0_4545 int_unitcell rval='r_int_cell' lval='l_int_cell' cval='c_int_cell'
xdint_5_1 ndint_x_909_4545 ndint_x_1818_4545 ndint_y_909_4545 ndint_y_909_5454 ndint_xy_909_4545 int_unitcell rval='r_int_cell' lval='l_int_cell' cval='c_int_cell'
xdint_5_2 ndint_x_1818_4545 ndint_x_2727_4545 ndint_y_1818_4545 ndint_y_1818_5454 ndint_xy_1818_4545 int_unitcell rval='r_int_cell' lval='l_int_cell' cval='c_int_cell'
xdint_5_3 ndint_x_2727_4545 ndint_x_3636_4545 ndint_y_2727_4545 ndint_y_2727_5454 ndint_xy_2727_4545 int_unitcell rval='r_int_cell' lval='l_int_cell' cval='c_int_cell'
xdint_5_4 ndint_x_3636_4545 ndint_x_4545_4545 ndint_y_3636_4545 ndint_y_3636_5454 ndint_xy_3636_4545 int_unitcell rval='r_int_cell' lval='l_int_cell' cval='c_int_cell'
xdint_5_5 ndint_x_4545_4545 ndint_x_5454_4545 ndint_y_4545_4545 ndint_y_4545_5454 ndint_xy_4545_4545 int_unitcell rval='r_int_cell' lval='l_int_cell' cval='c_int_cell'
xdint_5_6 ndint_x_5454_4545 ndint_x_6363_4545 ndint_y_5454_4545 ndint_y_5454_5454 ndint_xy_5454_4545 int_unitcell rval='r_int_cell' lval='l_int_cell' cval='c_int_cell'
xdint_5_7 ndint_x_6363_4545 ndint_x_7272_4545 ndint_y_6363_4545 ndint_y_6363_5454 ndint_xy_6363_4545 int_unitcell rval='r_int_cell' lval='l_int_cell' cval='c_int_cell'
xdint_5_8 ndint_x_7272_4545 ndint_x_8181_4545 ndint_y_7272_4545 ndint_y_7272_5454 ndint_xy_7272_4545 int_unitcell rval='r_int_cell' lval='l_int_cell' cval='c_int_cell'
xdint_5_9 ndint_x_8181_4545 ndint_x_9090_4545 ndint_y_8181_4545 ndint_y_8181_5454 ndint_xy_8181_4545 int_unitcell rval='r_int_cell' lval='l_int_cell' cval='c_int_cell'
xdint_5_10 ndint_x_9090_4545 ndint_x_9999_4545 ndint_y_9090_4545 ndint_y_9090_5454 ndint_xy_9090_4545 int_unitcell rval='r_int_cell' lval='l_int_cell' cval='c_int_cell'
xdint_6_0 ndint_x_0_5454 ndint_x_909_5454 ndint_y_0_5454 ndint_y_0_6363 ndint_xy_0_5454 int_unitcell rval='r_int_cell' lval='l_int_cell' cval='c_int_cell'
xdint_6_1 ndint_x_909_5454 ndint_x_1818_5454 ndint_y_909_5454 ndint_y_909_6363 ndint_xy_909_5454 int_unitcell rval='r_int_cell' lval='l_int_cell' cval='c_int_cell'
xdint_6_2 ndint_x_1818_5454 ndint_x_2727_5454 ndint_y_1818_5454 ndint_y_1818_6363 ndint_xy_1818_5454 int_unitcell rval='r_int_cell' lval='l_int_cell' cval='c_int_cell'
xdint_6_3 ndint_x_2727_5454 ndint_x_3636_5454 ndint_y_2727_5454 ndint_y_2727_6363 ndint_xy_2727_5454 int_unitcell rval='r_int_cell' lval='l_int_cell' cval='c_int_cell'
xdint_6_4 ndint_x_3636_5454 ndint_x_4545_5454 ndint_y_3636_5454 ndint_y_3636_6363 ndint_xy_3636_5454 int_unitcell rval='r_int_cell' lval='l_int_cell' cval='c_int_cell'
xdint_6_5 ndint_x_4545_5454 ndint_x_5454_5454 ndint_y_4545_5454 ndint_y_4545_6363 ndint_xy_4545_5454 int_unitcell rval='r_int_cell' lval='l_int_cell' cval='c_int_cell'
xdint_6_6 ndint_x_5454_5454 ndint_x_6363_5454 ndint_y_5454_5454 ndint_y_5454_6363 ndint_xy_5454_5454 int_unitcell rval='r_int_cell' lval='l_int_cell' cval='c_int_cell'
xdint_6_7 ndint_x_6363_5454 ndint_x_7272_5454 ndint_y_6363_5454 ndint_y_6363_6363 ndint_xy_6363_5454 int_unitcell rval='r_int_cell' lval='l_int_cell' cval='c_int_cell'
xdint_6_8 ndint_x_7272_5454 ndint_x_8181_5454 ndint_y_7272_5454 ndint_y_7272_6363 ndint_xy_7272_5454 int_unitcell rval='r_int_cell' lval='l_int_cell' cval='c_int_cell'
xdint_6_9 ndint_x_8181_5454 ndint_x_9090_5454 ndint_y_8181_5454 ndint_y_8181_6363 ndint_xy_8181_5454 int_unitcell rval='r_int_cell' lval='l_int_cell' cval='c_int_cell'
xdint_6_10 ndint_x_9090_5454 ndint_x_9999_5454 ndint_y_9090_5454 ndint_y_9090_6363 ndint_xy_9090_5454 int_unitcell rval='r_int_cell' lval='l_int_cell' cval='c_int_cell'
xdint_7_0 ndint_x_0_6363 ndint_x_909_6363 ndint_y_0_6363 ndint_y_0_7272 ndint_xy_0_6363 int_unitcell rval='r_int_cell' lval='l_int_cell' cval='c_int_cell'
xdint_7_1 ndint_x_909_6363 ndint_x_1818_6363 ndint_y_909_6363 ndint_y_909_7272 ndint_xy_909_6363 int_unitcell rval='r_int_cell' lval='l_int_cell' cval='c_int_cell'
xdint_7_2 ndint_x_1818_6363 ndint_x_2727_6363 ndint_y_1818_6363 ndint_y_1818_7272 ndint_xy_1818_6363 int_unitcell rval='r_int_cell' lval='l_int_cell' cval='c_int_cell'
xdint_7_3 ndint_x_2727_6363 ndint_x_3636_6363 ndint_y_2727_6363 ndint_y_2727_7272 ndint_xy_2727_6363 int_unitcell rval='r_int_cell' lval='l_int_cell' cval='c_int_cell'
xdint_7_4 ndint_x_3636_6363 ndint_x_4545_6363 ndint_y_3636_6363 ndint_y_3636_7272 ndint_xy_3636_6363 int_unitcell rval='r_int_cell' lval='l_int_cell' cval='c_int_cell'
xdint_7_5 ndint_x_4545_6363 ndint_x_5454_6363 ndint_y_4545_6363 ndint_y_4545_7272 ndint_xy_4545_6363 int_unitcell rval='r_int_cell' lval='l_int_cell' cval='c_int_cell'
xdint_7_6 ndint_x_5454_6363 ndint_x_6363_6363 ndint_y_5454_6363 ndint_y_5454_7272 ndint_xy_5454_6363 int_unitcell rval='r_int_cell' lval='l_int_cell' cval='c_int_cell'
xdint_7_7 ndint_x_6363_6363 ndint_x_7272_6363 ndint_y_6363_6363 ndint_y_6363_7272 ndint_xy_6363_6363 int_unitcell rval='r_int_cell' lval='l_int_cell' cval='c_int_cell'
xdint_7_8 ndint_x_7272_6363 ndint_x_8181_6363 ndint_y_7272_6363 ndint_y_7272_7272 ndint_xy_7272_6363 int_unitcell rval='r_int_cell' lval='l_int_cell' cval='c_int_cell'
xdint_7_9 ndint_x_8181_6363 ndint_x_9090_6363 ndint_y_8181_6363 ndint_y_8181_7272 ndint_xy_8181_6363 int_unitcell rval='r_int_cell' lval='l_int_cell' cval='c_int_cell'
xdint_7_10 ndint_x_9090_6363 ndint_x_9999_6363 ndint_y_9090_6363 ndint_y_9090_7272 ndint_xy_9090_6363 int_unitcell rval='r_int_cell' lval='l_int_cell' cval='c_int_cell'
xdint_8_0 ndint_x_0_7272 ndint_x_909_7272 ndint_y_0_7272 ndint_y_0_8181 ndint_xy_0_7272 int_unitcell rval='r_int_cell' lval='l_int_cell' cval='c_int_cell'
xdint_8_1 ndint_x_909_7272 ndint_x_1818_7272 ndint_y_909_7272 ndint_y_909_8181 ndint_xy_909_7272 int_unitcell rval='r_int_cell' lval='l_int_cell' cval='c_int_cell'
xdint_8_2 ndint_x_1818_7272 ndint_x_2727_7272 ndint_y_1818_7272 ndint_y_1818_8181 ndint_xy_1818_7272 int_unitcell rval='r_int_cell' lval='l_int_cell' cval='c_int_cell'
xdint_8_3 ndint_x_2727_7272 ndint_x_3636_7272 ndint_y_2727_7272 ndint_y_2727_8181 ndint_xy_2727_7272 int_unitcell rval='r_int_cell' lval='l_int_cell' cval='c_int_cell'
xdint_8_4 ndint_x_3636_7272 ndint_x_4545_7272 ndint_y_3636_7272 ndint_y_3636_8181 ndint_xy_3636_7272 int_unitcell rval='r_int_cell' lval='l_int_cell' cval='c_int_cell'
xdint_8_5 ndint_x_4545_7272 ndint_x_5454_7272 ndint_y_4545_7272 ndint_y_4545_8181 ndint_xy_4545_7272 int_unitcell rval='r_int_cell' lval='l_int_cell' cval='c_int_cell'
xdint_8_6 ndint_x_5454_7272 ndint_x_6363_7272 ndint_y_5454_7272 ndint_y_5454_8181 ndint_xy_5454_7272 int_unitcell rval='r_int_cell' lval='l_int_cell' cval='c_int_cell'
xdint_8_7 ndint_x_6363_7272 ndint_x_7272_7272 ndint_y_6363_7272 ndint_y_6363_8181 ndint_xy_6363_7272 int_unitcell rval='r_int_cell' lval='l_int_cell' cval='c_int_cell'
xdint_8_8 ndint_x_7272_7272 ndint_x_8181_7272 ndint_y_7272_7272 ndint_y_7272_8181 ndint_xy_7272_7272 int_unitcell rval='r_int_cell' lval='l_int_cell' cval='c_int_cell'
xdint_8_9 ndint_x_8181_7272 ndint_x_9090_7272 ndint_y_8181_7272 ndint_y_8181_8181 ndint_xy_8181_7272 int_unitcell rval='r_int_cell' lval='l_int_cell' cval='c_int_cell'
xdint_8_10 ndint_x_9090_7272 ndint_x_9999_7272 ndint_y_9090_7272 ndint_y_9090_8181 ndint_xy_9090_7272 int_unitcell rval='r_int_cell' lval='l_int_cell' cval='c_int_cell'
xdint_9_0 ndint_x_0_8181 ndint_x_909_8181 ndint_y_0_8181 ndint_y_0_9090 ndint_xy_0_8181 int_unitcell rval='r_int_cell' lval='l_int_cell' cval='c_int_cell'
xdint_9_1 ndint_x_909_8181 ndint_x_1818_8181 ndint_y_909_8181 ndint_y_909_9090 ndint_xy_909_8181 int_unitcell rval='r_int_cell' lval='l_int_cell' cval='c_int_cell'
xdint_9_2 ndint_x_1818_8181 ndint_x_2727_8181 ndint_y_1818_8181 ndint_y_1818_9090 ndint_xy_1818_8181 int_unitcell rval='r_int_cell' lval='l_int_cell' cval='c_int_cell'
xdint_9_3 ndint_x_2727_8181 ndint_x_3636_8181 ndint_y_2727_8181 ndint_y_2727_9090 ndint_xy_2727_8181 int_unitcell rval='r_int_cell' lval='l_int_cell' cval='c_int_cell'
xdint_9_4 ndint_x_3636_8181 ndint_x_4545_8181 ndint_y_3636_8181 ndint_y_3636_9090 ndint_xy_3636_8181 int_unitcell rval='r_int_cell' lval='l_int_cell' cval='c_int_cell'
xdint_9_5 ndint_x_4545_8181 ndint_x_5454_8181 ndint_y_4545_8181 ndint_y_4545_9090 ndint_xy_4545_8181 int_unitcell rval='r_int_cell' lval='l_int_cell' cval='c_int_cell'
xdint_9_6 ndint_x_5454_8181 ndint_x_6363_8181 ndint_y_5454_8181 ndint_y_5454_9090 ndint_xy_5454_8181 int_unitcell rval='r_int_cell' lval='l_int_cell' cval='c_int_cell'
xdint_9_7 ndint_x_6363_8181 ndint_x_7272_8181 ndint_y_6363_8181 ndint_y_6363_9090 ndint_xy_6363_8181 int_unitcell rval='r_int_cell' lval='l_int_cell' cval='c_int_cell'
xdint_9_8 ndint_x_7272_8181 ndint_x_8181_8181 ndint_y_7272_8181 ndint_y_7272_9090 ndint_xy_7272_8181 int_unitcell rval='r_int_cell' lval='l_int_cell' cval='c_int_cell'
xdint_9_9 ndint_x_8181_8181 ndint_x_9090_8181 ndint_y_8181_8181 ndint_y_8181_9090 ndint_xy_8181_8181 int_unitcell rval='r_int_cell' lval='l_int_cell' cval='c_int_cell'
xdint_9_10 ndint_x_9090_8181 ndint_x_9999_8181 ndint_y_9090_8181 ndint_y_9090_9090 ndint_xy_9090_8181 int_unitcell rval='r_int_cell' lval='l_int_cell' cval='c_int_cell'
xdint_10_0 ndint_x_0_9090 ndint_x_909_9090 ndint_y_0_9090 ndint_y_0_9999 ndint_xy_0_9090 int_unitcell rval='r_int_cell' lval='l_int_cell' cval='c_int_cell'
xdint_10_1 ndint_x_909_9090 ndint_x_1818_9090 ndint_y_909_9090 ndint_y_909_9999 ndint_xy_909_9090 int_unitcell rval='r_int_cell' lval='l_int_cell' cval='c_int_cell'
xdint_10_2 ndint_x_1818_9090 ndint_x_2727_9090 ndint_y_1818_9090 ndint_y_1818_9999 ndint_xy_1818_9090 int_unitcell rval='r_int_cell' lval='l_int_cell' cval='c_int_cell'
xdint_10_3 ndint_x_2727_9090 ndint_x_3636_9090 ndint_y_2727_9090 ndint_y_2727_9999 ndint_xy_2727_9090 int_unitcell rval='r_int_cell' lval='l_int_cell' cval='c_int_cell'
xdint_10_4 ndint_x_3636_9090 ndint_x_4545_9090 ndint_y_3636_9090 ndint_y_3636_9999 ndint_xy_3636_9090 int_unitcell rval='r_int_cell' lval='l_int_cell' cval='c_int_cell'
xdint_10_5 ndint_x_4545_9090 ndint_x_5454_9090 ndint_y_4545_9090 ndint_y_4545_9999 ndint_xy_4545_9090 int_unitcell rval='r_int_cell' lval='l_int_cell' cval='c_int_cell'
xdint_10_6 ndint_x_5454_9090 ndint_x_6363_9090 ndint_y_5454_9090 ndint_y_5454_9999 ndint_xy_5454_9090 int_unitcell rval='r_int_cell' lval='l_int_cell' cval='c_int_cell'
xdint_10_7 ndint_x_6363_9090 ndint_x_7272_9090 ndint_y_6363_9090 ndint_y_6363_9999 ndint_xy_6363_9090 int_unitcell rval='r_int_cell' lval='l_int_cell' cval='c_int_cell'
xdint_10_8 ndint_x_7272_9090 ndint_x_8181_9090 ndint_y_7272_9090 ndint_y_7272_9999 ndint_xy_7272_9090 int_unitcell rval='r_int_cell' lval='l_int_cell' cval='c_int_cell'
xdint_10_9 ndint_x_8181_9090 ndint_x_9090_9090 ndint_y_8181_9090 ndint_y_8181_9999 ndint_xy_8181_9090 int_unitcell rval='r_int_cell' lval='l_int_cell' cval='c_int_cell'
xdint_10_10 ndint_x_9090_9090 ndint_x_9999_9090 ndint_y_9090_9090 ndint_y_9090_9999 ndint_xy_9090_9090 int_unitcell rval='r_int_cell' lval='l_int_cell' cval='c_int_cell'


.include 'unitcell.subckt'

rd1_ubump2via_0_1 nd_chiplet1_pad_0_1 ndint_xy_909_909 0.001
rd1_ubump2via_0_3 nd_chiplet1_pad_0_3 ndint_y_909_1818 0.001
rd1_ubump2via_0_5 nd_chiplet1_pad_0_5 ndint_y_909_1818 0.001
rd1_ubump2via_0_7 nd_chiplet1_pad_0_7 ndint_y_909_1818 0.001
rd1_ubump2via_0_9 nd_chiplet1_pad_0_9 ndint_y_909_2727 0.001
rd1_ubump2via_1_0 nd_chiplet1_pad_1_0 ndint_y_1818_909 0.001
rd1_ubump2via_1_2 nd_chiplet1_pad_1_2 ndint_y_1818_1818 0.001
rd1_ubump2via_1_4 nd_chiplet1_pad_1_4 ndint_y_1818_1818 0.001
rd1_ubump2via_1_6 nd_chiplet1_pad_1_6 ndint_y_1818_1818 0.001
rd1_ubump2via_1_8 nd_chiplet1_pad_1_8 ndint_y_1818_2727 0.001
rd1_ubump2via_2_1 nd_chiplet1_pad_2_1 ndint_y_1818_909 0.001
rd1_ubump2via_2_3 nd_chiplet1_pad_2_3 ndint_y_1818_1818 0.001
rd1_ubump2via_2_5 nd_chiplet1_pad_2_5 ndint_xy_1818_1818 0.001
rd1_ubump2via_2_7 nd_chiplet1_pad_2_7 ndint_y_1818_1818 0.001
rd1_ubump2via_2_9 nd_chiplet1_pad_2_9 ndint_y_1818_2727 0.001
rd1_ubump2via_3_0 nd_chiplet1_pad_3_0 ndint_y_1818_909 0.001
rd1_ubump2via_3_2 nd_chiplet1_pad_3_2 ndint_y_1818_1818 0.001
rd1_ubump2via_3_4 nd_chiplet1_pad_3_4 ndint_y_1818_1818 0.001
rd1_ubump2via_3_6 nd_chiplet1_pad_3_6 ndint_y_1818_1818 0.001
rd1_ubump2via_3_8 nd_chiplet1_pad_3_8 ndint_y_1818_2727 0.001
rd1_ubump2via_4_1 nd_chiplet1_pad_4_1 ndint_y_2727_909 0.001
rd1_ubump2via_4_3 nd_chiplet1_pad_4_3 ndint_y_2727_1818 0.001
rd1_ubump2via_4_5 nd_chiplet1_pad_4_5 ndint_y_2727_1818 0.001
rd1_ubump2via_4_7 nd_chiplet1_pad_4_7 ndint_y_2727_1818 0.001
rd1_ubump2via_4_9 nd_chiplet1_pad_4_9 ndint_xy_2727_2727 0.001
rd1_ubump2via_5_0 nd_chiplet1_pad_5_0 ndint_xy_2727_909 0.001
rd1_ubump2via_5_2 nd_chiplet1_pad_5_2 ndint_y_2727_1818 0.001
rd1_ubump2via_5_4 nd_chiplet1_pad_5_4 ndint_y_2727_1818 0.001
rd1_ubump2via_5_6 nd_chiplet1_pad_5_6 ndint_y_2727_1818 0.001
rd1_ubump2via_5_8 nd_chiplet1_pad_5_8 ndint_y_2727_2727 0.001
rd1_ubump2via_6_1 nd_chiplet1_pad_6_1 ndint_y_3636_909 0.001
rd1_ubump2via_6_3 nd_chiplet1_pad_6_3 ndint_y_3636_1818 0.001
rd1_ubump2via_6_5 nd_chiplet1_pad_6_5 ndint_y_3636_1818 0.001
rd1_ubump2via_6_7 nd_chiplet1_pad_6_7 ndint_y_3636_1818 0.001
rd1_ubump2via_6_9 nd_chiplet1_pad_6_9 ndint_y_3636_2727 0.001
rd1_ubump2via_7_0 nd_chiplet1_pad_7_0 ndint_y_3636_909 0.001
rd1_ubump2via_7_2 nd_chiplet1_pad_7_2 ndint_y_3636_1818 0.001
rd1_ubump2via_7_4 nd_chiplet1_pad_7_4 ndint_xy_3636_1818 0.001
rd1_ubump2via_7_6 nd_chiplet1_pad_7_6 ndint_y_3636_1818 0.001
rd1_ubump2via_7_8 nd_chiplet1_pad_7_8 ndint_y_3636_2727 0.001
rd1_ubump2via_8_1 nd_chiplet1_pad_8_1 ndint_y_3636_909 0.001
rd1_ubump2via_8_3 nd_chiplet1_pad_8_3 ndint_y_3636_1818 0.001
rd1_ubump2via_8_5 nd_chiplet1_pad_8_5 ndint_y_3636_1818 0.001
rd1_ubump2via_8_7 nd_chiplet1_pad_8_7 ndint_y_3636_1818 0.001
rd1_ubump2via_8_9 nd_chiplet1_pad_8_9 ndint_y_3636_2727 0.001
rd1_ubump2via_9_0 nd_chiplet1_pad_9_0 ndint_y_4545_909 0.001
rd1_ubump2via_9_2 nd_chiplet1_pad_9_2 ndint_y_4545_1818 0.001
rd1_ubump2via_9_4 nd_chiplet1_pad_9_4 ndint_y_4545_1818 0.001
rd1_ubump2via_9_6 nd_chiplet1_pad_9_6 ndint_y_4545_1818 0.001
rd1_ubump2via_9_8 nd_chiplet1_pad_9_8 ndint_xy_4545_2727 0.001
rd2_ubump2via_0_1 nd_chiplet2_pad_0_1 ndint_xy_5454_909 0.001
rd2_ubump2via_0_3 nd_chiplet2_pad_0_3 ndint_y_5454_1818 0.001
rd2_ubump2via_0_5 nd_chiplet2_pad_0_5 ndint_y_5454_1818 0.001
rd2_ubump2via_0_7 nd_chiplet2_pad_0_7 ndint_y_5454_1818 0.001
rd2_ubump2via_0_9 nd_chiplet2_pad_0_9 ndint_y_5454_2727 0.001
rd2_ubump2via_1_0 nd_chiplet2_pad_1_0 ndint_y_6363_909 0.001
rd2_ubump2via_1_2 nd_chiplet2_pad_1_2 ndint_y_6363_1818 0.001
rd2_ubump2via_1_4 nd_chiplet2_pad_1_4 ndint_y_6363_1818 0.001
rd2_ubump2via_1_6 nd_chiplet2_pad_1_6 ndint_y_6363_1818 0.001
rd2_ubump2via_1_8 nd_chiplet2_pad_1_8 ndint_y_6363_2727 0.001
rd2_ubump2via_2_1 nd_chiplet2_pad_2_1 ndint_y_6363_909 0.001
rd2_ubump2via_2_3 nd_chiplet2_pad_2_3 ndint_y_6363_1818 0.001
rd2_ubump2via_2_5 nd_chiplet2_pad_2_5 ndint_xy_6363_1818 0.001
rd2_ubump2via_2_7 nd_chiplet2_pad_2_7 ndint_y_6363_1818 0.001
rd2_ubump2via_2_9 nd_chiplet2_pad_2_9 ndint_y_6363_2727 0.001
rd2_ubump2via_3_0 nd_chiplet2_pad_3_0 ndint_y_6363_909 0.001
rd2_ubump2via_3_2 nd_chiplet2_pad_3_2 ndint_y_6363_1818 0.001
rd2_ubump2via_3_4 nd_chiplet2_pad_3_4 ndint_y_6363_1818 0.001
rd2_ubump2via_3_6 nd_chiplet2_pad_3_6 ndint_y_6363_1818 0.001
rd2_ubump2via_3_8 nd_chiplet2_pad_3_8 ndint_y_6363_2727 0.001
rd2_ubump2via_4_1 nd_chiplet2_pad_4_1 ndint_y_7272_909 0.001
rd2_ubump2via_4_3 nd_chiplet2_pad_4_3 ndint_y_7272_1818 0.001
rd2_ubump2via_4_5 nd_chiplet2_pad_4_5 ndint_y_7272_1818 0.001
rd2_ubump2via_4_7 nd_chiplet2_pad_4_7 ndint_y_7272_1818 0.001
rd2_ubump2via_4_9 nd_chiplet2_pad_4_9 ndint_xy_7272_2727 0.001
rd2_ubump2via_5_0 nd_chiplet2_pad_5_0 ndint_xy_7272_909 0.001
rd2_ubump2via_5_2 nd_chiplet2_pad_5_2 ndint_y_7272_1818 0.001
rd2_ubump2via_5_4 nd_chiplet2_pad_5_4 ndint_y_7272_1818 0.001
rd2_ubump2via_5_6 nd_chiplet2_pad_5_6 ndint_y_7272_1818 0.001
rd2_ubump2via_5_8 nd_chiplet2_pad_5_8 ndint_y_7272_2727 0.001
rd2_ubump2via_6_1 nd_chiplet2_pad_6_1 ndint_y_8181_909 0.001
rd2_ubump2via_6_3 nd_chiplet2_pad_6_3 ndint_y_8181_1818 0.001
rd2_ubump2via_6_5 nd_chiplet2_pad_6_5 ndint_y_8181_1818 0.001
rd2_ubump2via_6_7 nd_chiplet2_pad_6_7 ndint_y_8181_1818 0.001
rd2_ubump2via_6_9 nd_chiplet2_pad_6_9 ndint_y_8181_2727 0.001
rd2_ubump2via_7_0 nd_chiplet2_pad_7_0 ndint_y_8181_909 0.001
rd2_ubump2via_7_2 nd_chiplet2_pad_7_2 ndint_y_8181_1818 0.001
rd2_ubump2via_7_4 nd_chiplet2_pad_7_4 ndint_xy_8181_1818 0.001
rd2_ubump2via_7_6 nd_chiplet2_pad_7_6 ndint_y_8181_1818 0.001
rd2_ubump2via_7_8 nd_chiplet2_pad_7_8 ndint_y_8181_2727 0.001
rd2_ubump2via_8_1 nd_chiplet2_pad_8_1 ndint_y_8181_909 0.001
rd2_ubump2via_8_3 nd_chiplet2_pad_8_3 ndint_y_8181_1818 0.001
rd2_ubump2via_8_5 nd_chiplet2_pad_8_5 ndint_y_8181_1818 0.001
rd2_ubump2via_8_7 nd_chiplet2_pad_8_7 ndint_y_8181_1818 0.001
rd2_ubump2via_8_9 nd_chiplet2_pad_8_9 ndint_y_8181_2727 0.001
rd2_ubump2via_9_0 nd_chiplet2_pad_9_0 ndint_y_9090_909 0.001
rd2_ubump2via_9_2 nd_chiplet2_pad_9_2 ndint_y_9090_1818 0.001
rd2_ubump2via_9_4 nd_chiplet2_pad_9_4 ndint_y_9090_1818 0.001
rd2_ubump2via_9_6 nd_chiplet2_pad_9_6 ndint_y_9090_1818 0.001
rd2_ubump2via_9_8 nd_chiplet2_pad_9_8 ndint_xy_9090_2727 0.001
rd3_ubump2via_0_1 nd_chiplet3_pad_0_1 ndint_y_1818_4545 0.001
rd3_ubump2via_0_3 nd_chiplet3_pad_0_3 ndint_y_1818_4545 0.001
rd3_ubump2via_0_5 nd_chiplet3_pad_0_5 ndint_y_1818_5454 0.001
rd3_ubump2via_0_7 nd_chiplet3_pad_0_7 ndint_y_1818_5454 0.001
rd3_ubump2via_0_9 nd_chiplet3_pad_0_9 ndint_y_1818_6363 0.001
rd3_ubump2via_1_0 nd_chiplet3_pad_1_0 ndint_y_2727_3636 0.001
rd3_ubump2via_1_2 nd_chiplet3_pad_1_2 ndint_y_2727_4545 0.001
rd3_ubump2via_1_4 nd_chiplet3_pad_1_4 ndint_y_2727_4545 0.001
rd3_ubump2via_1_6 nd_chiplet3_pad_1_6 ndint_y_2727_5454 0.001
rd3_ubump2via_1_8 nd_chiplet3_pad_1_8 ndint_y_2727_5454 0.001
rd3_ubump2via_2_1 nd_chiplet3_pad_2_1 ndint_y_2727_4545 0.001
rd3_ubump2via_2_3 nd_chiplet3_pad_2_3 ndint_y_2727_4545 0.001
rd3_ubump2via_2_5 nd_chiplet3_pad_2_5 ndint_y_2727_5454 0.001
rd3_ubump2via_2_7 nd_chiplet3_pad_2_7 ndint_y_2727_5454 0.001
rd3_ubump2via_2_9 nd_chiplet3_pad_2_9 ndint_y_2727_6363 0.001
rd3_ubump2via_3_0 nd_chiplet3_pad_3_0 ndint_y_2727_3636 0.001
rd3_ubump2via_3_2 nd_chiplet3_pad_3_2 ndint_y_2727_4545 0.001
rd3_ubump2via_3_4 nd_chiplet3_pad_3_4 ndint_y_2727_4545 0.001
rd3_ubump2via_3_6 nd_chiplet3_pad_3_6 ndint_y_2727_5454 0.001
rd3_ubump2via_3_8 nd_chiplet3_pad_3_8 ndint_y_2727_5454 0.001
rd3_ubump2via_4_1 nd_chiplet3_pad_4_1 ndint_y_2727_4545 0.001
rd3_ubump2via_4_3 nd_chiplet3_pad_4_3 ndint_y_2727_4545 0.001
rd3_ubump2via_4_5 nd_chiplet3_pad_4_5 ndint_y_2727_5454 0.001
rd3_ubump2via_4_7 nd_chiplet3_pad_4_7 ndint_y_2727_5454 0.001
rd3_ubump2via_4_9 nd_chiplet3_pad_4_9 ndint_y_2727_6363 0.001
rd3_ubump2via_5_0 nd_chiplet3_pad_5_0 ndint_y_3636_3636 0.001
rd3_ubump2via_5_2 nd_chiplet3_pad_5_2 ndint_y_3636_4545 0.001
rd3_ubump2via_5_4 nd_chiplet3_pad_5_4 ndint_y_3636_4545 0.001
rd3_ubump2via_5_6 nd_chiplet3_pad_5_6 ndint_y_3636_5454 0.001
rd3_ubump2via_5_8 nd_chiplet3_pad_5_8 ndint_y_3636_5454 0.001
rd3_ubump2via_6_1 nd_chiplet3_pad_6_1 ndint_y_3636_4545 0.001
rd3_ubump2via_6_3 nd_chiplet3_pad_6_3 ndint_y_3636_4545 0.001
rd3_ubump2via_6_5 nd_chiplet3_pad_6_5 ndint_y_3636_5454 0.001
rd3_ubump2via_6_7 nd_chiplet3_pad_6_7 ndint_y_3636_5454 0.001
rd3_ubump2via_6_9 nd_chiplet3_pad_6_9 ndint_y_3636_6363 0.001
rd3_ubump2via_7_0 nd_chiplet3_pad_7_0 ndint_y_3636_3636 0.001
rd3_ubump2via_7_2 nd_chiplet3_pad_7_2 ndint_y_3636_4545 0.001
rd3_ubump2via_7_4 nd_chiplet3_pad_7_4 ndint_y_3636_4545 0.001
rd3_ubump2via_7_6 nd_chiplet3_pad_7_6 ndint_y_3636_5454 0.001
rd3_ubump2via_7_8 nd_chiplet3_pad_7_8 ndint_y_3636_5454 0.001
rd3_ubump2via_8_1 nd_chiplet3_pad_8_1 ndint_y_3636_4545 0.001
rd3_ubump2via_8_3 nd_chiplet3_pad_8_3 ndint_y_3636_4545 0.001
rd3_ubump2via_8_5 nd_chiplet3_pad_8_5 ndint_y_3636_5454 0.001
rd3_ubump2via_8_7 nd_chiplet3_pad_8_7 ndint_y_3636_5454 0.001
rd3_ubump2via_8_9 nd_chiplet3_pad_8_9 ndint_y_3636_6363 0.001
rd3_ubump2via_9_0 nd_chiplet3_pad_9_0 ndint_y_4545_3636 0.001
rd3_ubump2via_9_2 nd_chiplet3_pad_9_2 ndint_y_4545_4545 0.001
rd3_ubump2via_9_4 nd_chiplet3_pad_9_4 ndint_y_4545_4545 0.001
rd3_ubump2via_9_6 nd_chiplet3_pad_9_6 ndint_y_4545_5454 0.001
rd3_ubump2via_9_8 nd_chiplet3_pad_9_8 ndint_y_4545_5454 0.001
rd4_ubump2via_0_1 nd_chiplet4_pad_0_1 ndint_y_5454_4545 0.001
rd4_ubump2via_0_3 nd_chiplet4_pad_0_3 ndint_y_5454_4545 0.001
rd4_ubump2via_0_5 nd_chiplet4_pad_0_5 ndint_y_5454_5454 0.001
rd4_ubump2via_0_7 nd_chiplet4_pad_0_7 ndint_y_5454_5454 0.001
rd4_ubump2via_0_9 nd_chiplet4_pad_0_9 ndint_y_5454_6363 0.001
rd4_ubump2via_1_0 nd_chiplet4_pad_1_0 ndint_y_6363_3636 0.001
rd4_ubump2via_1_2 nd_chiplet4_pad_1_2 ndint_y_6363_4545 0.001
rd4_ubump2via_1_4 nd_chiplet4_pad_1_4 ndint_y_6363_4545 0.001
rd4_ubump2via_1_6 nd_chiplet4_pad_1_6 ndint_y_6363_5454 0.001
rd4_ubump2via_1_8 nd_chiplet4_pad_1_8 ndint_y_6363_5454 0.001
rd4_ubump2via_2_1 nd_chiplet4_pad_2_1 ndint_y_6363_4545 0.001
rd4_ubump2via_2_3 nd_chiplet4_pad_2_3 ndint_y_6363_4545 0.001
rd4_ubump2via_2_5 nd_chiplet4_pad_2_5 ndint_y_6363_5454 0.001
rd4_ubump2via_2_7 nd_chiplet4_pad_2_7 ndint_y_6363_5454 0.001
rd4_ubump2via_2_9 nd_chiplet4_pad_2_9 ndint_y_6363_6363 0.001
rd4_ubump2via_3_0 nd_chiplet4_pad_3_0 ndint_y_6363_3636 0.001
rd4_ubump2via_3_2 nd_chiplet4_pad_3_2 ndint_y_6363_4545 0.001
rd4_ubump2via_3_4 nd_chiplet4_pad_3_4 ndint_y_6363_4545 0.001
rd4_ubump2via_3_6 nd_chiplet4_pad_3_6 ndint_y_6363_5454 0.001
rd4_ubump2via_3_8 nd_chiplet4_pad_3_8 ndint_y_6363_5454 0.001
rd4_ubump2via_4_1 nd_chiplet4_pad_4_1 ndint_y_6363_4545 0.001
rd4_ubump2via_4_3 nd_chiplet4_pad_4_3 ndint_y_6363_4545 0.001
rd4_ubump2via_4_5 nd_chiplet4_pad_4_5 ndint_y_6363_5454 0.001
rd4_ubump2via_4_7 nd_chiplet4_pad_4_7 ndint_y_6363_5454 0.001
rd4_ubump2via_4_9 nd_chiplet4_pad_4_9 ndint_y_6363_6363 0.001
rd4_ubump2via_5_0 nd_chiplet4_pad_5_0 ndint_y_7272_3636 0.001
rd4_ubump2via_5_2 nd_chiplet4_pad_5_2 ndint_y_7272_4545 0.001
rd4_ubump2via_5_4 nd_chiplet4_pad_5_4 ndint_y_7272_4545 0.001
rd4_ubump2via_5_6 nd_chiplet4_pad_5_6 ndint_y_7272_5454 0.001
rd4_ubump2via_5_8 nd_chiplet4_pad_5_8 ndint_y_7272_5454 0.001
rd4_ubump2via_6_1 nd_chiplet4_pad_6_1 ndint_y_7272_4545 0.001
rd4_ubump2via_6_3 nd_chiplet4_pad_6_3 ndint_y_7272_4545 0.001
rd4_ubump2via_6_5 nd_chiplet4_pad_6_5 ndint_y_7272_5454 0.001
rd4_ubump2via_6_7 nd_chiplet4_pad_6_7 ndint_y_7272_5454 0.001
rd4_ubump2via_6_9 nd_chiplet4_pad_6_9 ndint_y_7272_6363 0.001
rd4_ubump2via_7_0 nd_chiplet4_pad_7_0 ndint_y_7272_3636 0.001
rd4_ubump2via_7_2 nd_chiplet4_pad_7_2 ndint_y_7272_4545 0.001
rd4_ubump2via_7_4 nd_chiplet4_pad_7_4 ndint_y_7272_4545 0.001
rd4_ubump2via_7_6 nd_chiplet4_pad_7_6 ndint_y_7272_5454 0.001
rd4_ubump2via_7_8 nd_chiplet4_pad_7_8 ndint_y_7272_5454 0.001
rd4_ubump2via_8_1 nd_chiplet4_pad_8_1 ndint_y_7272_4545 0.001
rd4_ubump2via_8_3 nd_chiplet4_pad_8_3 ndint_y_7272_4545 0.001
rd4_ubump2via_8_5 nd_chiplet4_pad_8_5 ndint_y_7272_5454 0.001
rd4_ubump2via_8_7 nd_chiplet4_pad_8_7 ndint_y_7272_5454 0.001
rd4_ubump2via_8_9 nd_chiplet4_pad_8_9 ndint_y_7272_6363 0.001
rd4_ubump2via_9_0 nd_chiplet4_pad_9_0 ndint_y_8181_3636 0.001
rd4_ubump2via_9_2 nd_chiplet4_pad_9_2 ndint_y_8181_4545 0.001
rd4_ubump2via_9_4 nd_chiplet4_pad_9_4 ndint_y_8181_4545 0.001
rd4_ubump2via_9_6 nd_chiplet4_pad_9_6 ndint_y_8181_5454 0.001
rd4_ubump2via_9_8 nd_chiplet4_pad_9_8 ndint_y_8181_5454 0.001
rd5_ubump2via_0_1 nd_chiplet5_pad_0_1 ndint_xy_909_7272 0.001
rd5_ubump2via_0_3 nd_chiplet5_pad_0_3 ndint_y_909_8181 0.001
rd5_ubump2via_0_5 nd_chiplet5_pad_0_5 ndint_y_909_8181 0.001
rd5_ubump2via_0_7 nd_chiplet5_pad_0_7 ndint_y_909_8181 0.001
rd5_ubump2via_0_9 nd_chiplet5_pad_0_9 ndint_y_909_9090 0.001
rd5_ubump2via_1_0 nd_chiplet5_pad_1_0 ndint_y_1818_7272 0.001
rd5_ubump2via_1_2 nd_chiplet5_pad_1_2 ndint_y_1818_8181 0.001
rd5_ubump2via_1_4 nd_chiplet5_pad_1_4 ndint_y_1818_8181 0.001
rd5_ubump2via_1_6 nd_chiplet5_pad_1_6 ndint_y_1818_8181 0.001
rd5_ubump2via_1_8 nd_chiplet5_pad_1_8 ndint_y_1818_9090 0.001
rd5_ubump2via_2_1 nd_chiplet5_pad_2_1 ndint_y_1818_7272 0.001
rd5_ubump2via_2_3 nd_chiplet5_pad_2_3 ndint_y_1818_8181 0.001
rd5_ubump2via_2_5 nd_chiplet5_pad_2_5 ndint_xy_1818_8181 0.001
rd5_ubump2via_2_7 nd_chiplet5_pad_2_7 ndint_y_1818_8181 0.001
rd5_ubump2via_2_9 nd_chiplet5_pad_2_9 ndint_y_1818_9090 0.001
rd5_ubump2via_3_0 nd_chiplet5_pad_3_0 ndint_y_1818_7272 0.001
rd5_ubump2via_3_2 nd_chiplet5_pad_3_2 ndint_y_1818_8181 0.001
rd5_ubump2via_3_4 nd_chiplet5_pad_3_4 ndint_y_1818_8181 0.001
rd5_ubump2via_3_6 nd_chiplet5_pad_3_6 ndint_y_1818_8181 0.001
rd5_ubump2via_3_8 nd_chiplet5_pad_3_8 ndint_y_1818_9090 0.001
rd5_ubump2via_4_1 nd_chiplet5_pad_4_1 ndint_y_2727_7272 0.001
rd5_ubump2via_4_3 nd_chiplet5_pad_4_3 ndint_y_2727_8181 0.001
rd5_ubump2via_4_5 nd_chiplet5_pad_4_5 ndint_y_2727_8181 0.001
rd5_ubump2via_4_7 nd_chiplet5_pad_4_7 ndint_y_2727_8181 0.001
rd5_ubump2via_4_9 nd_chiplet5_pad_4_9 ndint_xy_2727_9090 0.001
rd5_ubump2via_5_0 nd_chiplet5_pad_5_0 ndint_xy_2727_7272 0.001
rd5_ubump2via_5_2 nd_chiplet5_pad_5_2 ndint_y_2727_8181 0.001
rd5_ubump2via_5_4 nd_chiplet5_pad_5_4 ndint_y_2727_8181 0.001
rd5_ubump2via_5_6 nd_chiplet5_pad_5_6 ndint_y_2727_8181 0.001
rd5_ubump2via_5_8 nd_chiplet5_pad_5_8 ndint_y_2727_9090 0.001
rd5_ubump2via_6_1 nd_chiplet5_pad_6_1 ndint_y_3636_7272 0.001
rd5_ubump2via_6_3 nd_chiplet5_pad_6_3 ndint_y_3636_8181 0.001
rd5_ubump2via_6_5 nd_chiplet5_pad_6_5 ndint_y_3636_8181 0.001
rd5_ubump2via_6_7 nd_chiplet5_pad_6_7 ndint_y_3636_8181 0.001
rd5_ubump2via_6_9 nd_chiplet5_pad_6_9 ndint_y_3636_9090 0.001
rd5_ubump2via_7_0 nd_chiplet5_pad_7_0 ndint_y_3636_7272 0.001
rd5_ubump2via_7_2 nd_chiplet5_pad_7_2 ndint_y_3636_8181 0.001
rd5_ubump2via_7_4 nd_chiplet5_pad_7_4 ndint_xy_3636_8181 0.001
rd5_ubump2via_7_6 nd_chiplet5_pad_7_6 ndint_y_3636_8181 0.001
rd5_ubump2via_7_8 nd_chiplet5_pad_7_8 ndint_y_3636_9090 0.001
rd5_ubump2via_8_1 nd_chiplet5_pad_8_1 ndint_y_3636_7272 0.001
rd5_ubump2via_8_3 nd_chiplet5_pad_8_3 ndint_y_3636_8181 0.001
rd5_ubump2via_8_5 nd_chiplet5_pad_8_5 ndint_y_3636_8181 0.001
rd5_ubump2via_8_7 nd_chiplet5_pad_8_7 ndint_y_3636_8181 0.001
rd5_ubump2via_8_9 nd_chiplet5_pad_8_9 ndint_y_3636_9090 0.001
rd5_ubump2via_9_0 nd_chiplet5_pad_9_0 ndint_y_4545_7272 0.001
rd5_ubump2via_9_2 nd_chiplet5_pad_9_2 ndint_y_4545_8181 0.001
rd5_ubump2via_9_4 nd_chiplet5_pad_9_4 ndint_y_4545_8181 0.001
rd5_ubump2via_9_6 nd_chiplet5_pad_9_6 ndint_y_4545_8181 0.001
rd5_ubump2via_9_8 nd_chiplet5_pad_9_8 ndint_xy_4545_9090 0.001
rd6_ubump2via_0_1 nd_chiplet6_pad_0_1 ndint_xy_5454_7272 0.001
rd6_ubump2via_0_3 nd_chiplet6_pad_0_3 ndint_y_5454_8181 0.001
rd6_ubump2via_0_5 nd_chiplet6_pad_0_5 ndint_y_5454_8181 0.001
rd6_ubump2via_0_7 nd_chiplet6_pad_0_7 ndint_y_5454_8181 0.001
rd6_ubump2via_0_9 nd_chiplet6_pad_0_9 ndint_y_5454_9090 0.001
rd6_ubump2via_1_0 nd_chiplet6_pad_1_0 ndint_y_6363_7272 0.001
rd6_ubump2via_1_2 nd_chiplet6_pad_1_2 ndint_y_6363_8181 0.001
rd6_ubump2via_1_4 nd_chiplet6_pad_1_4 ndint_y_6363_8181 0.001
rd6_ubump2via_1_6 nd_chiplet6_pad_1_6 ndint_y_6363_8181 0.001
rd6_ubump2via_1_8 nd_chiplet6_pad_1_8 ndint_y_6363_9090 0.001
rd6_ubump2via_2_1 nd_chiplet6_pad_2_1 ndint_y_6363_7272 0.001
rd6_ubump2via_2_3 nd_chiplet6_pad_2_3 ndint_y_6363_8181 0.001
rd6_ubump2via_2_5 nd_chiplet6_pad_2_5 ndint_xy_6363_8181 0.001
rd6_ubump2via_2_7 nd_chiplet6_pad_2_7 ndint_y_6363_8181 0.001
rd6_ubump2via_2_9 nd_chiplet6_pad_2_9 ndint_y_6363_9090 0.001
rd6_ubump2via_3_0 nd_chiplet6_pad_3_0 ndint_y_6363_7272 0.001
rd6_ubump2via_3_2 nd_chiplet6_pad_3_2 ndint_y_6363_8181 0.001
rd6_ubump2via_3_4 nd_chiplet6_pad_3_4 ndint_y_6363_8181 0.001
rd6_ubump2via_3_6 nd_chiplet6_pad_3_6 ndint_y_6363_8181 0.001
rd6_ubump2via_3_8 nd_chiplet6_pad_3_8 ndint_y_6363_9090 0.001
rd6_ubump2via_4_1 nd_chiplet6_pad_4_1 ndint_y_7272_7272 0.001
rd6_ubump2via_4_3 nd_chiplet6_pad_4_3 ndint_y_7272_8181 0.001
rd6_ubump2via_4_5 nd_chiplet6_pad_4_5 ndint_y_7272_8181 0.001
rd6_ubump2via_4_7 nd_chiplet6_pad_4_7 ndint_y_7272_8181 0.001
rd6_ubump2via_4_9 nd_chiplet6_pad_4_9 ndint_xy_7272_9090 0.001
rd6_ubump2via_5_0 nd_chiplet6_pad_5_0 ndint_xy_7272_7272 0.001
rd6_ubump2via_5_2 nd_chiplet6_pad_5_2 ndint_y_7272_8181 0.001
rd6_ubump2via_5_4 nd_chiplet6_pad_5_4 ndint_y_7272_8181 0.001
rd6_ubump2via_5_6 nd_chiplet6_pad_5_6 ndint_y_7272_8181 0.001
rd6_ubump2via_5_8 nd_chiplet6_pad_5_8 ndint_y_7272_9090 0.001
rd6_ubump2via_6_1 nd_chiplet6_pad_6_1 ndint_y_8181_7272 0.001
rd6_ubump2via_6_3 nd_chiplet6_pad_6_3 ndint_y_8181_8181 0.001
rd6_ubump2via_6_5 nd_chiplet6_pad_6_5 ndint_y_8181_8181 0.001
rd6_ubump2via_6_7 nd_chiplet6_pad_6_7 ndint_y_8181_8181 0.001
rd6_ubump2via_6_9 nd_chiplet6_pad_6_9 ndint_y_8181_9090 0.001
rd6_ubump2via_7_0 nd_chiplet6_pad_7_0 ndint_y_8181_7272 0.001
rd6_ubump2via_7_2 nd_chiplet6_pad_7_2 ndint_y_8181_8181 0.001
rd6_ubump2via_7_4 nd_chiplet6_pad_7_4 ndint_xy_8181_8181 0.001
rd6_ubump2via_7_6 nd_chiplet6_pad_7_6 ndint_y_8181_8181 0.001
rd6_ubump2via_7_8 nd_chiplet6_pad_7_8 ndint_y_8181_9090 0.001
rd6_ubump2via_8_1 nd_chiplet6_pad_8_1 ndint_y_8181_7272 0.001
rd6_ubump2via_8_3 nd_chiplet6_pad_8_3 ndint_y_8181_8181 0.001
rd6_ubump2via_8_5 nd_chiplet6_pad_8_5 ndint_y_8181_8181 0.001
rd6_ubump2via_8_7 nd_chiplet6_pad_8_7 ndint_y_8181_8181 0.001
rd6_ubump2via_8_9 nd_chiplet6_pad_8_9 ndint_y_8181_9090 0.001
rd6_ubump2via_9_0 nd_chiplet6_pad_9_0 ndint_y_9090_7272 0.001
rd6_ubump2via_9_2 nd_chiplet6_pad_9_2 ndint_y_9090_8181 0.001
rd6_ubump2via_9_4 nd_chiplet6_pad_9_4 ndint_y_9090_8181 0.001
rd6_ubump2via_9_6 nd_chiplet6_pad_9_6 ndint_y_9090_8181 0.001
rd6_ubump2via_9_8 nd_chiplet6_pad_9_8 ndint_xy_9090_9090 0.001

*-- chiplet instance [0]: chiplet1
xchiplet_chiplet1
+nd_chiplet1_pad_0_1
+nd_chiplet1_pad_0_3
+nd_chiplet1_pad_0_5
+nd_chiplet1_pad_0_7
+nd_chiplet1_pad_0_9
+nd_chiplet1_pad_1_0
+nd_chiplet1_pad_1_2
+nd_chiplet1_pad_1_4
+nd_chiplet1_pad_1_6
+nd_chiplet1_pad_1_8
+nd_chiplet1_pad_2_1
+nd_chiplet1_pad_2_3
+nd_chiplet1_pad_2_5
+nd_chiplet1_pad_2_7
+nd_chiplet1_pad_2_9
+nd_chiplet1_pad_3_0
+nd_chiplet1_pad_3_2
+nd_chiplet1_pad_3_4
+nd_chiplet1_pad_3_6
+nd_chiplet1_pad_3_8
+nd_chiplet1_pad_4_1
+nd_chiplet1_pad_4_3
+nd_chiplet1_pad_4_5
+nd_chiplet1_pad_4_7
+nd_chiplet1_pad_4_9
+nd_chiplet1_pad_5_0
+nd_chiplet1_pad_5_2
+nd_chiplet1_pad_5_4
+nd_chiplet1_pad_5_6
+nd_chiplet1_pad_5_8
+nd_chiplet1_pad_6_1
+nd_chiplet1_pad_6_3
+nd_chiplet1_pad_6_5
+nd_chiplet1_pad_6_7
+nd_chiplet1_pad_6_9
+nd_chiplet1_pad_7_0
+nd_chiplet1_pad_7_2
+nd_chiplet1_pad_7_4
+nd_chiplet1_pad_7_6
+nd_chiplet1_pad_7_8
+nd_chiplet1_pad_8_1
+nd_chiplet1_pad_8_3
+nd_chiplet1_pad_8_5
+nd_chiplet1_pad_8_7
+nd_chiplet1_pad_8_9
+nd_chiplet1_pad_9_0
+nd_chiplet1_pad_9_2
+nd_chiplet1_pad_9_4
+nd_chiplet1_pad_9_6
+nd_chiplet1_pad_9_8
+chiplet1

*-- chiplet instance [1]: chiplet2
xchiplet_chiplet2
+nd_chiplet2_pad_0_1
+nd_chiplet2_pad_0_3
+nd_chiplet2_pad_0_5
+nd_chiplet2_pad_0_7
+nd_chiplet2_pad_0_9
+nd_chiplet2_pad_1_0
+nd_chiplet2_pad_1_2
+nd_chiplet2_pad_1_4
+nd_chiplet2_pad_1_6
+nd_chiplet2_pad_1_8
+nd_chiplet2_pad_2_1
+nd_chiplet2_pad_2_3
+nd_chiplet2_pad_2_5
+nd_chiplet2_pad_2_7
+nd_chiplet2_pad_2_9
+nd_chiplet2_pad_3_0
+nd_chiplet2_pad_3_2
+nd_chiplet2_pad_3_4
+nd_chiplet2_pad_3_6
+nd_chiplet2_pad_3_8
+nd_chiplet2_pad_4_1
+nd_chiplet2_pad_4_3
+nd_chiplet2_pad_4_5
+nd_chiplet2_pad_4_7
+nd_chiplet2_pad_4_9
+nd_chiplet2_pad_5_0
+nd_chiplet2_pad_5_2
+nd_chiplet2_pad_5_4
+nd_chiplet2_pad_5_6
+nd_chiplet2_pad_5_8
+nd_chiplet2_pad_6_1
+nd_chiplet2_pad_6_3
+nd_chiplet2_pad_6_5
+nd_chiplet2_pad_6_7
+nd_chiplet2_pad_6_9
+nd_chiplet2_pad_7_0
+nd_chiplet2_pad_7_2
+nd_chiplet2_pad_7_4
+nd_chiplet2_pad_7_6
+nd_chiplet2_pad_7_8
+nd_chiplet2_pad_8_1
+nd_chiplet2_pad_8_3
+nd_chiplet2_pad_8_5
+nd_chiplet2_pad_8_7
+nd_chiplet2_pad_8_9
+nd_chiplet2_pad_9_0
+nd_chiplet2_pad_9_2
+nd_chiplet2_pad_9_4
+nd_chiplet2_pad_9_6
+nd_chiplet2_pad_9_8
+chiplet2

*-- chiplet instance [2]: chiplet3
xchiplet_chiplet3
+nd_chiplet3_pad_0_1
+nd_chiplet3_pad_0_3
+nd_chiplet3_pad_0_5
+nd_chiplet3_pad_0_7
+nd_chiplet3_pad_0_9
+nd_chiplet3_pad_1_0
+nd_chiplet3_pad_1_2
+nd_chiplet3_pad_1_4
+nd_chiplet3_pad_1_6
+nd_chiplet3_pad_1_8
+nd_chiplet3_pad_2_1
+nd_chiplet3_pad_2_3
+nd_chiplet3_pad_2_5
+nd_chiplet3_pad_2_7
+nd_chiplet3_pad_2_9
+nd_chiplet3_pad_3_0
+nd_chiplet3_pad_3_2
+nd_chiplet3_pad_3_4
+nd_chiplet3_pad_3_6
+nd_chiplet3_pad_3_8
+nd_chiplet3_pad_4_1
+nd_chiplet3_pad_4_3
+nd_chiplet3_pad_4_5
+nd_chiplet3_pad_4_7
+nd_chiplet3_pad_4_9
+nd_chiplet3_pad_5_0
+nd_chiplet3_pad_5_2
+nd_chiplet3_pad_5_4
+nd_chiplet3_pad_5_6
+nd_chiplet3_pad_5_8
+nd_chiplet3_pad_6_1
+nd_chiplet3_pad_6_3
+nd_chiplet3_pad_6_5
+nd_chiplet3_pad_6_7
+nd_chiplet3_pad_6_9
+nd_chiplet3_pad_7_0
+nd_chiplet3_pad_7_2
+nd_chiplet3_pad_7_4
+nd_chiplet3_pad_7_6
+nd_chiplet3_pad_7_8
+nd_chiplet3_pad_8_1
+nd_chiplet3_pad_8_3
+nd_chiplet3_pad_8_5
+nd_chiplet3_pad_8_7
+nd_chiplet3_pad_8_9
+nd_chiplet3_pad_9_0
+nd_chiplet3_pad_9_2
+nd_chiplet3_pad_9_4
+nd_chiplet3_pad_9_6
+nd_chiplet3_pad_9_8
+chiplet3

*-- chiplet instance [3]: chiplet4
xchiplet_chiplet4
+nd_chiplet4_pad_0_1
+nd_chiplet4_pad_0_3
+nd_chiplet4_pad_0_5
+nd_chiplet4_pad_0_7
+nd_chiplet4_pad_0_9
+nd_chiplet4_pad_1_0
+nd_chiplet4_pad_1_2
+nd_chiplet4_pad_1_4
+nd_chiplet4_pad_1_6
+nd_chiplet4_pad_1_8
+nd_chiplet4_pad_2_1
+nd_chiplet4_pad_2_3
+nd_chiplet4_pad_2_5
+nd_chiplet4_pad_2_7
+nd_chiplet4_pad_2_9
+nd_chiplet4_pad_3_0
+nd_chiplet4_pad_3_2
+nd_chiplet4_pad_3_4
+nd_chiplet4_pad_3_6
+nd_chiplet4_pad_3_8
+nd_chiplet4_pad_4_1
+nd_chiplet4_pad_4_3
+nd_chiplet4_pad_4_5
+nd_chiplet4_pad_4_7
+nd_chiplet4_pad_4_9
+nd_chiplet4_pad_5_0
+nd_chiplet4_pad_5_2
+nd_chiplet4_pad_5_4
+nd_chiplet4_pad_5_6
+nd_chiplet4_pad_5_8
+nd_chiplet4_pad_6_1
+nd_chiplet4_pad_6_3
+nd_chiplet4_pad_6_5
+nd_chiplet4_pad_6_7
+nd_chiplet4_pad_6_9
+nd_chiplet4_pad_7_0
+nd_chiplet4_pad_7_2
+nd_chiplet4_pad_7_4
+nd_chiplet4_pad_7_6
+nd_chiplet4_pad_7_8
+nd_chiplet4_pad_8_1
+nd_chiplet4_pad_8_3
+nd_chiplet4_pad_8_5
+nd_chiplet4_pad_8_7
+nd_chiplet4_pad_8_9
+nd_chiplet4_pad_9_0
+nd_chiplet4_pad_9_2
+nd_chiplet4_pad_9_4
+nd_chiplet4_pad_9_6
+nd_chiplet4_pad_9_8
+chiplet4

*-- chiplet instance [4]: chiplet5
xchiplet_chiplet5
+nd_chiplet5_pad_0_1
+nd_chiplet5_pad_0_3
+nd_chiplet5_pad_0_5
+nd_chiplet5_pad_0_7
+nd_chiplet5_pad_0_9
+nd_chiplet5_pad_1_0
+nd_chiplet5_pad_1_2
+nd_chiplet5_pad_1_4
+nd_chiplet5_pad_1_6
+nd_chiplet5_pad_1_8
+nd_chiplet5_pad_2_1
+nd_chiplet5_pad_2_3
+nd_chiplet5_pad_2_5
+nd_chiplet5_pad_2_7
+nd_chiplet5_pad_2_9
+nd_chiplet5_pad_3_0
+nd_chiplet5_pad_3_2
+nd_chiplet5_pad_3_4
+nd_chiplet5_pad_3_6
+nd_chiplet5_pad_3_8
+nd_chiplet5_pad_4_1
+nd_chiplet5_pad_4_3
+nd_chiplet5_pad_4_5
+nd_chiplet5_pad_4_7
+nd_chiplet5_pad_4_9
+nd_chiplet5_pad_5_0
+nd_chiplet5_pad_5_2
+nd_chiplet5_pad_5_4
+nd_chiplet5_pad_5_6
+nd_chiplet5_pad_5_8
+nd_chiplet5_pad_6_1
+nd_chiplet5_pad_6_3
+nd_chiplet5_pad_6_5
+nd_chiplet5_pad_6_7
+nd_chiplet5_pad_6_9
+nd_chiplet5_pad_7_0
+nd_chiplet5_pad_7_2
+nd_chiplet5_pad_7_4
+nd_chiplet5_pad_7_6
+nd_chiplet5_pad_7_8
+nd_chiplet5_pad_8_1
+nd_chiplet5_pad_8_3
+nd_chiplet5_pad_8_5
+nd_chiplet5_pad_8_7
+nd_chiplet5_pad_8_9
+nd_chiplet5_pad_9_0
+nd_chiplet5_pad_9_2
+nd_chiplet5_pad_9_4
+nd_chiplet5_pad_9_6
+nd_chiplet5_pad_9_8
+chiplet5

*-- chiplet instance [5]: chiplet6
xchiplet_chiplet6
+nd_chiplet6_pad_0_1
+nd_chiplet6_pad_0_3
+nd_chiplet6_pad_0_5
+nd_chiplet6_pad_0_7
+nd_chiplet6_pad_0_9
+nd_chiplet6_pad_1_0
+nd_chiplet6_pad_1_2
+nd_chiplet6_pad_1_4
+nd_chiplet6_pad_1_6
+nd_chiplet6_pad_1_8
+nd_chiplet6_pad_2_1
+nd_chiplet6_pad_2_3
+nd_chiplet6_pad_2_5
+nd_chiplet6_pad_2_7
+nd_chiplet6_pad_2_9
+nd_chiplet6_pad_3_0
+nd_chiplet6_pad_3_2
+nd_chiplet6_pad_3_4
+nd_chiplet6_pad_3_6
+nd_chiplet6_pad_3_8
+nd_chiplet6_pad_4_1
+nd_chiplet6_pad_4_3
+nd_chiplet6_pad_4_5
+nd_chiplet6_pad_4_7
+nd_chiplet6_pad_4_9
+nd_chiplet6_pad_5_0
+nd_chiplet6_pad_5_2
+nd_chiplet6_pad_5_4
+nd_chiplet6_pad_5_6
+nd_chiplet6_pad_5_8
+nd_chiplet6_pad_6_1
+nd_chiplet6_pad_6_3
+nd_chiplet6_pad_6_5
+nd_chiplet6_pad_6_7
+nd_chiplet6_pad_6_9
+nd_chiplet6_pad_7_0
+nd_chiplet6_pad_7_2
+nd_chiplet6_pad_7_4
+nd_chiplet6_pad_7_6
+nd_chiplet6_pad_7_8
+nd_chiplet6_pad_8_1
+nd_chiplet6_pad_8_3
+nd_chiplet6_pad_8_5
+nd_chiplet6_pad_8_7
+nd_chiplet6_pad_8_9
+nd_chiplet6_pad_9_0
+nd_chiplet6_pad_9_2
+nd_chiplet6_pad_9_4
+nd_chiplet6_pad_9_6
+nd_chiplet6_pad_9_8
+chiplet6
.include 'chiplet1_ac.subckt'
.include 'chiplet2_ac.subckt'
.include 'chiplet3_ac.subckt'
.include 'chiplet4_ac.subckt'
.include 'chiplet5_ac.subckt'
.include 'chiplet6_ac.subckt'

*-- tsv array
xdint_tsv_0_1 ndint_tsv_0_1 ndint_bump_0_1 int_tsv
xdint_tsv_0_3 ndint_tsv_0_3 ndint_bump_0_3 int_tsv
xdint_tsv_0_5 ndint_tsv_0_5 ndint_bump_0_5 int_tsv
xdint_tsv_0_7 ndint_tsv_0_7 ndint_bump_0_7 int_tsv
xdint_tsv_0_9 ndint_tsv_0_9 ndint_bump_0_9 int_tsv
xdint_tsv_0_11 ndint_tsv_0_11 ndint_bump_0_11 int_tsv
xdint_tsv_0_13 ndint_tsv_0_13 ndint_bump_0_13 int_tsv
xdint_tsv_0_15 ndint_tsv_0_15 ndint_bump_0_15 int_tsv
xdint_tsv_0_17 ndint_tsv_0_17 ndint_bump_0_17 int_tsv
xdint_tsv_0_19 ndint_tsv_0_19 ndint_bump_0_19 int_tsv
xdint_tsv_1_0 ndint_tsv_1_0 ndint_bump_1_0 int_tsv
xdint_tsv_1_2 ndint_tsv_1_2 ndint_bump_1_2 int_tsv
xdint_tsv_1_4 ndint_tsv_1_4 ndint_bump_1_4 int_tsv
xdint_tsv_1_6 ndint_tsv_1_6 ndint_bump_1_6 int_tsv
xdint_tsv_1_8 ndint_tsv_1_8 ndint_bump_1_8 int_tsv
xdint_tsv_1_10 ndint_tsv_1_10 ndint_bump_1_10 int_tsv
xdint_tsv_1_12 ndint_tsv_1_12 ndint_bump_1_12 int_tsv
xdint_tsv_1_14 ndint_tsv_1_14 ndint_bump_1_14 int_tsv
xdint_tsv_1_16 ndint_tsv_1_16 ndint_bump_1_16 int_tsv
xdint_tsv_1_18 ndint_tsv_1_18 ndint_bump_1_18 int_tsv
xdint_tsv_2_1 ndint_tsv_2_1 ndint_bump_2_1 int_tsv
xdint_tsv_2_3 ndint_tsv_2_3 ndint_bump_2_3 int_tsv
xdint_tsv_2_5 ndint_tsv_2_5 ndint_bump_2_5 int_tsv
xdint_tsv_2_7 ndint_tsv_2_7 ndint_bump_2_7 int_tsv
xdint_tsv_2_9 ndint_tsv_2_9 ndint_bump_2_9 int_tsv
xdint_tsv_2_11 ndint_tsv_2_11 ndint_bump_2_11 int_tsv
xdint_tsv_2_13 ndint_tsv_2_13 ndint_bump_2_13 int_tsv
xdint_tsv_2_15 ndint_tsv_2_15 ndint_bump_2_15 int_tsv
xdint_tsv_2_17 ndint_tsv_2_17 ndint_bump_2_17 int_tsv
xdint_tsv_2_19 ndint_tsv_2_19 ndint_bump_2_19 int_tsv
xdint_tsv_3_0 ndint_tsv_3_0 ndint_bump_3_0 int_tsv
xdint_tsv_3_2 ndint_tsv_3_2 ndint_bump_3_2 int_tsv
xdint_tsv_3_4 ndint_tsv_3_4 ndint_bump_3_4 int_tsv
xdint_tsv_3_6 ndint_tsv_3_6 ndint_bump_3_6 int_tsv
xdint_tsv_3_8 ndint_tsv_3_8 ndint_bump_3_8 int_tsv
xdint_tsv_3_10 ndint_tsv_3_10 ndint_bump_3_10 int_tsv
xdint_tsv_3_12 ndint_tsv_3_12 ndint_bump_3_12 int_tsv
xdint_tsv_3_14 ndint_tsv_3_14 ndint_bump_3_14 int_tsv
xdint_tsv_3_16 ndint_tsv_3_16 ndint_bump_3_16 int_tsv
xdint_tsv_3_18 ndint_tsv_3_18 ndint_bump_3_18 int_tsv
xdint_tsv_4_1 ndint_tsv_4_1 ndint_bump_4_1 int_tsv
xdint_tsv_4_3 ndint_tsv_4_3 ndint_bump_4_3 int_tsv
xdint_tsv_4_5 ndint_tsv_4_5 ndint_bump_4_5 int_tsv
xdint_tsv_4_7 ndint_tsv_4_7 ndint_bump_4_7 int_tsv
xdint_tsv_4_9 ndint_tsv_4_9 ndint_bump_4_9 int_tsv
xdint_tsv_4_11 ndint_tsv_4_11 ndint_bump_4_11 int_tsv
xdint_tsv_4_13 ndint_tsv_4_13 ndint_bump_4_13 int_tsv
xdint_tsv_4_15 ndint_tsv_4_15 ndint_bump_4_15 int_tsv
xdint_tsv_4_17 ndint_tsv_4_17 ndint_bump_4_17 int_tsv
xdint_tsv_4_19 ndint_tsv_4_19 ndint_bump_4_19 int_tsv
xdint_tsv_5_0 ndint_tsv_5_0 ndint_bump_5_0 int_tsv
xdint_tsv_5_2 ndint_tsv_5_2 ndint_bump_5_2 int_tsv
xdint_tsv_5_4 ndint_tsv_5_4 ndint_bump_5_4 int_tsv
xdint_tsv_5_6 ndint_tsv_5_6 ndint_bump_5_6 int_tsv
xdint_tsv_5_8 ndint_tsv_5_8 ndint_bump_5_8 int_tsv
xdint_tsv_5_10 ndint_tsv_5_10 ndint_bump_5_10 int_tsv
xdint_tsv_5_12 ndint_tsv_5_12 ndint_bump_5_12 int_tsv
xdint_tsv_5_14 ndint_tsv_5_14 ndint_bump_5_14 int_tsv
xdint_tsv_5_16 ndint_tsv_5_16 ndint_bump_5_16 int_tsv
xdint_tsv_5_18 ndint_tsv_5_18 ndint_bump_5_18 int_tsv
xdint_tsv_6_1 ndint_tsv_6_1 ndint_bump_6_1 int_tsv
xdint_tsv_6_3 ndint_tsv_6_3 ndint_bump_6_3 int_tsv
xdint_tsv_6_5 ndint_tsv_6_5 ndint_bump_6_5 int_tsv
xdint_tsv_6_7 ndint_tsv_6_7 ndint_bump_6_7 int_tsv
xdint_tsv_6_9 ndint_tsv_6_9 ndint_bump_6_9 int_tsv
xdint_tsv_6_11 ndint_tsv_6_11 ndint_bump_6_11 int_tsv
xdint_tsv_6_13 ndint_tsv_6_13 ndint_bump_6_13 int_tsv
xdint_tsv_6_15 ndint_tsv_6_15 ndint_bump_6_15 int_tsv
xdint_tsv_6_17 ndint_tsv_6_17 ndint_bump_6_17 int_tsv
xdint_tsv_6_19 ndint_tsv_6_19 ndint_bump_6_19 int_tsv
xdint_tsv_7_0 ndint_tsv_7_0 ndint_bump_7_0 int_tsv
xdint_tsv_7_2 ndint_tsv_7_2 ndint_bump_7_2 int_tsv
xdint_tsv_7_4 ndint_tsv_7_4 ndint_bump_7_4 int_tsv
xdint_tsv_7_6 ndint_tsv_7_6 ndint_bump_7_6 int_tsv
xdint_tsv_7_8 ndint_tsv_7_8 ndint_bump_7_8 int_tsv
xdint_tsv_7_10 ndint_tsv_7_10 ndint_bump_7_10 int_tsv
xdint_tsv_7_12 ndint_tsv_7_12 ndint_bump_7_12 int_tsv
xdint_tsv_7_14 ndint_tsv_7_14 ndint_bump_7_14 int_tsv
xdint_tsv_7_16 ndint_tsv_7_16 ndint_bump_7_16 int_tsv
xdint_tsv_7_18 ndint_tsv_7_18 ndint_bump_7_18 int_tsv
xdint_tsv_8_1 ndint_tsv_8_1 ndint_bump_8_1 int_tsv
xdint_tsv_8_3 ndint_tsv_8_3 ndint_bump_8_3 int_tsv
xdint_tsv_8_5 ndint_tsv_8_5 ndint_bump_8_5 int_tsv
xdint_tsv_8_7 ndint_tsv_8_7 ndint_bump_8_7 int_tsv
xdint_tsv_8_9 ndint_tsv_8_9 ndint_bump_8_9 int_tsv
xdint_tsv_8_11 ndint_tsv_8_11 ndint_bump_8_11 int_tsv
xdint_tsv_8_13 ndint_tsv_8_13 ndint_bump_8_13 int_tsv
xdint_tsv_8_15 ndint_tsv_8_15 ndint_bump_8_15 int_tsv
xdint_tsv_8_17 ndint_tsv_8_17 ndint_bump_8_17 int_tsv
xdint_tsv_8_19 ndint_tsv_8_19 ndint_bump_8_19 int_tsv
xdint_tsv_9_0 ndint_tsv_9_0 ndint_bump_9_0 int_tsv
xdint_tsv_9_2 ndint_tsv_9_2 ndint_bump_9_2 int_tsv
xdint_tsv_9_4 ndint_tsv_9_4 ndint_bump_9_4 int_tsv
xdint_tsv_9_6 ndint_tsv_9_6 ndint_bump_9_6 int_tsv
xdint_tsv_9_8 ndint_tsv_9_8 ndint_bump_9_8 int_tsv
xdint_tsv_9_10 ndint_tsv_9_10 ndint_bump_9_10 int_tsv
xdint_tsv_9_12 ndint_tsv_9_12 ndint_bump_9_12 int_tsv
xdint_tsv_9_14 ndint_tsv_9_14 ndint_bump_9_14 int_tsv
xdint_tsv_9_16 ndint_tsv_9_16 ndint_bump_9_16 int_tsv
xdint_tsv_9_18 ndint_tsv_9_18 ndint_bump_9_18 int_tsv
xdint_tsv_10_1 ndint_tsv_10_1 ndint_bump_10_1 int_tsv
xdint_tsv_10_3 ndint_tsv_10_3 ndint_bump_10_3 int_tsv
xdint_tsv_10_5 ndint_tsv_10_5 ndint_bump_10_5 int_tsv
xdint_tsv_10_7 ndint_tsv_10_7 ndint_bump_10_7 int_tsv
xdint_tsv_10_9 ndint_tsv_10_9 ndint_bump_10_9 int_tsv
xdint_tsv_10_11 ndint_tsv_10_11 ndint_bump_10_11 int_tsv
xdint_tsv_10_13 ndint_tsv_10_13 ndint_bump_10_13 int_tsv
xdint_tsv_10_15 ndint_tsv_10_15 ndint_bump_10_15 int_tsv
xdint_tsv_10_17 ndint_tsv_10_17 ndint_bump_10_17 int_tsv
xdint_tsv_10_19 ndint_tsv_10_19 ndint_bump_10_19 int_tsv
xdint_tsv_11_0 ndint_tsv_11_0 ndint_bump_11_0 int_tsv
xdint_tsv_11_2 ndint_tsv_11_2 ndint_bump_11_2 int_tsv
xdint_tsv_11_4 ndint_tsv_11_4 ndint_bump_11_4 int_tsv
xdint_tsv_11_6 ndint_tsv_11_6 ndint_bump_11_6 int_tsv
xdint_tsv_11_8 ndint_tsv_11_8 ndint_bump_11_8 int_tsv
xdint_tsv_11_10 ndint_tsv_11_10 ndint_bump_11_10 int_tsv
xdint_tsv_11_12 ndint_tsv_11_12 ndint_bump_11_12 int_tsv
xdint_tsv_11_14 ndint_tsv_11_14 ndint_bump_11_14 int_tsv
xdint_tsv_11_16 ndint_tsv_11_16 ndint_bump_11_16 int_tsv
xdint_tsv_11_18 ndint_tsv_11_18 ndint_bump_11_18 int_tsv
xdint_tsv_12_1 ndint_tsv_12_1 ndint_bump_12_1 int_tsv
xdint_tsv_12_3 ndint_tsv_12_3 ndint_bump_12_3 int_tsv
xdint_tsv_12_5 ndint_tsv_12_5 ndint_bump_12_5 int_tsv
xdint_tsv_12_7 ndint_tsv_12_7 ndint_bump_12_7 int_tsv
xdint_tsv_12_9 ndint_tsv_12_9 ndint_bump_12_9 int_tsv
xdint_tsv_12_11 ndint_tsv_12_11 ndint_bump_12_11 int_tsv
xdint_tsv_12_13 ndint_tsv_12_13 ndint_bump_12_13 int_tsv
xdint_tsv_12_15 ndint_tsv_12_15 ndint_bump_12_15 int_tsv
xdint_tsv_12_17 ndint_tsv_12_17 ndint_bump_12_17 int_tsv
xdint_tsv_12_19 ndint_tsv_12_19 ndint_bump_12_19 int_tsv
xdint_tsv_13_0 ndint_tsv_13_0 ndint_bump_13_0 int_tsv
xdint_tsv_13_2 ndint_tsv_13_2 ndint_bump_13_2 int_tsv
xdint_tsv_13_4 ndint_tsv_13_4 ndint_bump_13_4 int_tsv
xdint_tsv_13_6 ndint_tsv_13_6 ndint_bump_13_6 int_tsv
xdint_tsv_13_8 ndint_tsv_13_8 ndint_bump_13_8 int_tsv
xdint_tsv_13_10 ndint_tsv_13_10 ndint_bump_13_10 int_tsv
xdint_tsv_13_12 ndint_tsv_13_12 ndint_bump_13_12 int_tsv
xdint_tsv_13_14 ndint_tsv_13_14 ndint_bump_13_14 int_tsv
xdint_tsv_13_16 ndint_tsv_13_16 ndint_bump_13_16 int_tsv
xdint_tsv_13_18 ndint_tsv_13_18 ndint_bump_13_18 int_tsv
xdint_tsv_14_1 ndint_tsv_14_1 ndint_bump_14_1 int_tsv
xdint_tsv_14_3 ndint_tsv_14_3 ndint_bump_14_3 int_tsv
xdint_tsv_14_5 ndint_tsv_14_5 ndint_bump_14_5 int_tsv
xdint_tsv_14_7 ndint_tsv_14_7 ndint_bump_14_7 int_tsv
xdint_tsv_14_9 ndint_tsv_14_9 ndint_bump_14_9 int_tsv
xdint_tsv_14_11 ndint_tsv_14_11 ndint_bump_14_11 int_tsv
xdint_tsv_14_13 ndint_tsv_14_13 ndint_bump_14_13 int_tsv
xdint_tsv_14_15 ndint_tsv_14_15 ndint_bump_14_15 int_tsv
xdint_tsv_14_17 ndint_tsv_14_17 ndint_bump_14_17 int_tsv
xdint_tsv_14_19 ndint_tsv_14_19 ndint_bump_14_19 int_tsv
xdint_tsv_15_0 ndint_tsv_15_0 ndint_bump_15_0 int_tsv
xdint_tsv_15_2 ndint_tsv_15_2 ndint_bump_15_2 int_tsv
xdint_tsv_15_4 ndint_tsv_15_4 ndint_bump_15_4 int_tsv
xdint_tsv_15_6 ndint_tsv_15_6 ndint_bump_15_6 int_tsv
xdint_tsv_15_8 ndint_tsv_15_8 ndint_bump_15_8 int_tsv
xdint_tsv_15_10 ndint_tsv_15_10 ndint_bump_15_10 int_tsv
xdint_tsv_15_12 ndint_tsv_15_12 ndint_bump_15_12 int_tsv
xdint_tsv_15_14 ndint_tsv_15_14 ndint_bump_15_14 int_tsv
xdint_tsv_15_16 ndint_tsv_15_16 ndint_bump_15_16 int_tsv
xdint_tsv_15_18 ndint_tsv_15_18 ndint_bump_15_18 int_tsv
xdint_tsv_16_1 ndint_tsv_16_1 ndint_bump_16_1 int_tsv
xdint_tsv_16_3 ndint_tsv_16_3 ndint_bump_16_3 int_tsv
xdint_tsv_16_5 ndint_tsv_16_5 ndint_bump_16_5 int_tsv
xdint_tsv_16_7 ndint_tsv_16_7 ndint_bump_16_7 int_tsv
xdint_tsv_16_9 ndint_tsv_16_9 ndint_bump_16_9 int_tsv
xdint_tsv_16_11 ndint_tsv_16_11 ndint_bump_16_11 int_tsv
xdint_tsv_16_13 ndint_tsv_16_13 ndint_bump_16_13 int_tsv
xdint_tsv_16_15 ndint_tsv_16_15 ndint_bump_16_15 int_tsv
xdint_tsv_16_17 ndint_tsv_16_17 ndint_bump_16_17 int_tsv
xdint_tsv_16_19 ndint_tsv_16_19 ndint_bump_16_19 int_tsv
xdint_tsv_17_0 ndint_tsv_17_0 ndint_bump_17_0 int_tsv
xdint_tsv_17_2 ndint_tsv_17_2 ndint_bump_17_2 int_tsv
xdint_tsv_17_4 ndint_tsv_17_4 ndint_bump_17_4 int_tsv
xdint_tsv_17_6 ndint_tsv_17_6 ndint_bump_17_6 int_tsv
xdint_tsv_17_8 ndint_tsv_17_8 ndint_bump_17_8 int_tsv
xdint_tsv_17_10 ndint_tsv_17_10 ndint_bump_17_10 int_tsv
xdint_tsv_17_12 ndint_tsv_17_12 ndint_bump_17_12 int_tsv
xdint_tsv_17_14 ndint_tsv_17_14 ndint_bump_17_14 int_tsv
xdint_tsv_17_16 ndint_tsv_17_16 ndint_bump_17_16 int_tsv
xdint_tsv_17_18 ndint_tsv_17_18 ndint_bump_17_18 int_tsv
xdint_tsv_18_1 ndint_tsv_18_1 ndint_bump_18_1 int_tsv
xdint_tsv_18_3 ndint_tsv_18_3 ndint_bump_18_3 int_tsv
xdint_tsv_18_5 ndint_tsv_18_5 ndint_bump_18_5 int_tsv
xdint_tsv_18_7 ndint_tsv_18_7 ndint_bump_18_7 int_tsv
xdint_tsv_18_9 ndint_tsv_18_9 ndint_bump_18_9 int_tsv
xdint_tsv_18_11 ndint_tsv_18_11 ndint_bump_18_11 int_tsv
xdint_tsv_18_13 ndint_tsv_18_13 ndint_bump_18_13 int_tsv
xdint_tsv_18_15 ndint_tsv_18_15 ndint_bump_18_15 int_tsv
xdint_tsv_18_17 ndint_tsv_18_17 ndint_bump_18_17 int_tsv
xdint_tsv_18_19 ndint_tsv_18_19 ndint_bump_18_19 int_tsv
xdint_tsv_19_0 ndint_tsv_19_0 ndint_bump_19_0 int_tsv
xdint_tsv_19_2 ndint_tsv_19_2 ndint_bump_19_2 int_tsv
xdint_tsv_19_4 ndint_tsv_19_4 ndint_bump_19_4 int_tsv
xdint_tsv_19_6 ndint_tsv_19_6 ndint_bump_19_6 int_tsv
xdint_tsv_19_8 ndint_tsv_19_8 ndint_bump_19_8 int_tsv
xdint_tsv_19_10 ndint_tsv_19_10 ndint_bump_19_10 int_tsv
xdint_tsv_19_12 ndint_tsv_19_12 ndint_bump_19_12 int_tsv
xdint_tsv_19_14 ndint_tsv_19_14 ndint_bump_19_14 int_tsv
xdint_tsv_19_16 ndint_tsv_19_16 ndint_bump_19_16 int_tsv
xdint_tsv_19_18 ndint_tsv_19_18 ndint_bump_19_18 int_tsv
.include 'int_tsv.subckt'

*-- tsv to via
rdint_tsv2via_0_1 ndint_tsv_0_1 ndint_y_909_909 0.001
rdint_tsv2via_0_3 ndint_tsv_0_3 ndint_y_909_1818 0.001
rdint_tsv2via_0_5 ndint_tsv_0_5 ndint_y_909_2727 0.001
rdint_tsv2via_0_7 ndint_tsv_0_7 ndint_y_909_3636 0.001
rdint_tsv2via_0_9 ndint_tsv_0_9 ndint_y_909_4545 0.001
rdint_tsv2via_0_11 ndint_tsv_0_11 ndint_y_909_5454 0.001
rdint_tsv2via_0_13 ndint_tsv_0_13 ndint_y_909_6363 0.001
rdint_tsv2via_0_15 ndint_tsv_0_15 ndint_y_909_7272 0.001
rdint_tsv2via_0_17 ndint_tsv_0_17 ndint_y_909_8181 0.001
rdint_tsv2via_0_19 ndint_tsv_0_19 ndint_xy_909_9090 0.001
rdint_tsv2via_1_0 ndint_tsv_1_0 ndint_y_909_909 0.001
rdint_tsv2via_1_2 ndint_tsv_1_2 ndint_y_909_1818 0.001
rdint_tsv2via_1_4 ndint_tsv_1_4 ndint_y_909_2727 0.001
rdint_tsv2via_1_6 ndint_tsv_1_6 ndint_y_909_3636 0.001
rdint_tsv2via_1_8 ndint_tsv_1_8 ndint_y_909_4545 0.001
rdint_tsv2via_1_10 ndint_tsv_1_10 ndint_y_909_5454 0.001
rdint_tsv2via_1_12 ndint_tsv_1_12 ndint_y_909_6363 0.001
rdint_tsv2via_1_14 ndint_tsv_1_14 ndint_y_909_7272 0.001
rdint_tsv2via_1_16 ndint_tsv_1_16 ndint_y_909_8181 0.001
rdint_tsv2via_1_18 ndint_tsv_1_18 ndint_xy_909_9090 0.001
rdint_tsv2via_2_1 ndint_tsv_2_1 ndint_y_1818_909 0.001
rdint_tsv2via_2_3 ndint_tsv_2_3 ndint_y_1818_1818 0.001
rdint_tsv2via_2_5 ndint_tsv_2_5 ndint_y_1818_2727 0.001
rdint_tsv2via_2_7 ndint_tsv_2_7 ndint_y_1818_3636 0.001
rdint_tsv2via_2_9 ndint_tsv_2_9 ndint_y_1818_4545 0.001
rdint_tsv2via_2_11 ndint_tsv_2_11 ndint_y_1818_5454 0.001
rdint_tsv2via_2_13 ndint_tsv_2_13 ndint_y_1818_6363 0.001
rdint_tsv2via_2_15 ndint_tsv_2_15 ndint_y_1818_7272 0.001
rdint_tsv2via_2_17 ndint_tsv_2_17 ndint_xy_1818_8181 0.001
rdint_tsv2via_2_19 ndint_tsv_2_19 ndint_y_1818_9090 0.001
rdint_tsv2via_3_0 ndint_tsv_3_0 ndint_y_1818_909 0.001
rdint_tsv2via_3_2 ndint_tsv_3_2 ndint_y_1818_1818 0.001
rdint_tsv2via_3_4 ndint_tsv_3_4 ndint_y_1818_2727 0.001
rdint_tsv2via_3_6 ndint_tsv_3_6 ndint_y_1818_3636 0.001
rdint_tsv2via_3_8 ndint_tsv_3_8 ndint_y_1818_4545 0.001
rdint_tsv2via_3_10 ndint_tsv_3_10 ndint_y_1818_5454 0.001
rdint_tsv2via_3_12 ndint_tsv_3_12 ndint_y_1818_6363 0.001
rdint_tsv2via_3_14 ndint_tsv_3_14 ndint_y_1818_7272 0.001
rdint_tsv2via_3_16 ndint_tsv_3_16 ndint_xy_1818_8181 0.001
rdint_tsv2via_3_18 ndint_tsv_3_18 ndint_y_1818_9090 0.001
rdint_tsv2via_4_1 ndint_tsv_4_1 ndint_y_2727_909 0.001
rdint_tsv2via_4_3 ndint_tsv_4_3 ndint_y_2727_1818 0.001
rdint_tsv2via_4_5 ndint_tsv_4_5 ndint_y_2727_2727 0.001
rdint_tsv2via_4_7 ndint_tsv_4_7 ndint_y_2727_3636 0.001
rdint_tsv2via_4_9 ndint_tsv_4_9 ndint_y_2727_4545 0.001
rdint_tsv2via_4_11 ndint_tsv_4_11 ndint_y_2727_5454 0.001
rdint_tsv2via_4_13 ndint_tsv_4_13 ndint_y_2727_6363 0.001
rdint_tsv2via_4_15 ndint_tsv_4_15 ndint_xy_2727_7272 0.001
rdint_tsv2via_4_17 ndint_tsv_4_17 ndint_y_2727_8181 0.001
rdint_tsv2via_4_19 ndint_tsv_4_19 ndint_y_2727_9090 0.001
rdint_tsv2via_5_0 ndint_tsv_5_0 ndint_y_2727_909 0.001
rdint_tsv2via_5_2 ndint_tsv_5_2 ndint_y_2727_1818 0.001
rdint_tsv2via_5_4 ndint_tsv_5_4 ndint_y_2727_2727 0.001
rdint_tsv2via_5_6 ndint_tsv_5_6 ndint_y_2727_3636 0.001
rdint_tsv2via_5_8 ndint_tsv_5_8 ndint_y_2727_4545 0.001
rdint_tsv2via_5_10 ndint_tsv_5_10 ndint_y_2727_5454 0.001
rdint_tsv2via_5_12 ndint_tsv_5_12 ndint_y_2727_6363 0.001
rdint_tsv2via_5_14 ndint_tsv_5_14 ndint_xy_2727_7272 0.001
rdint_tsv2via_5_16 ndint_tsv_5_16 ndint_y_2727_8181 0.001
rdint_tsv2via_5_18 ndint_tsv_5_18 ndint_y_2727_9090 0.001
rdint_tsv2via_6_1 ndint_tsv_6_1 ndint_y_3636_909 0.001
rdint_tsv2via_6_3 ndint_tsv_6_3 ndint_y_3636_1818 0.001
rdint_tsv2via_6_5 ndint_tsv_6_5 ndint_y_3636_2727 0.001
rdint_tsv2via_6_7 ndint_tsv_6_7 ndint_y_3636_3636 0.001
rdint_tsv2via_6_9 ndint_tsv_6_9 ndint_y_3636_4545 0.001
rdint_tsv2via_6_11 ndint_tsv_6_11 ndint_y_3636_5454 0.001
rdint_tsv2via_6_13 ndint_tsv_6_13 ndint_xy_3636_6363 0.001
rdint_tsv2via_6_15 ndint_tsv_6_15 ndint_y_3636_7272 0.001
rdint_tsv2via_6_17 ndint_tsv_6_17 ndint_y_3636_8181 0.001
rdint_tsv2via_6_19 ndint_tsv_6_19 ndint_y_3636_9090 0.001
rdint_tsv2via_7_0 ndint_tsv_7_0 ndint_y_3636_909 0.001
rdint_tsv2via_7_2 ndint_tsv_7_2 ndint_y_3636_1818 0.001
rdint_tsv2via_7_4 ndint_tsv_7_4 ndint_y_3636_2727 0.001
rdint_tsv2via_7_6 ndint_tsv_7_6 ndint_y_3636_3636 0.001
rdint_tsv2via_7_8 ndint_tsv_7_8 ndint_y_3636_4545 0.001
rdint_tsv2via_7_10 ndint_tsv_7_10 ndint_y_3636_5454 0.001
rdint_tsv2via_7_12 ndint_tsv_7_12 ndint_xy_3636_6363 0.001
rdint_tsv2via_7_14 ndint_tsv_7_14 ndint_y_3636_7272 0.001
rdint_tsv2via_7_16 ndint_tsv_7_16 ndint_y_3636_8181 0.001
rdint_tsv2via_7_18 ndint_tsv_7_18 ndint_y_3636_9090 0.001
rdint_tsv2via_8_1 ndint_tsv_8_1 ndint_y_4545_909 0.001
rdint_tsv2via_8_3 ndint_tsv_8_3 ndint_y_4545_1818 0.001
rdint_tsv2via_8_5 ndint_tsv_8_5 ndint_y_4545_2727 0.001
rdint_tsv2via_8_7 ndint_tsv_8_7 ndint_y_4545_3636 0.001
rdint_tsv2via_8_9 ndint_tsv_8_9 ndint_y_4545_4545 0.001
rdint_tsv2via_8_11 ndint_tsv_8_11 ndint_xy_4545_5454 0.001
rdint_tsv2via_8_13 ndint_tsv_8_13 ndint_y_4545_6363 0.001
rdint_tsv2via_8_15 ndint_tsv_8_15 ndint_y_4545_7272 0.001
rdint_tsv2via_8_17 ndint_tsv_8_17 ndint_y_4545_8181 0.001
rdint_tsv2via_8_19 ndint_tsv_8_19 ndint_y_4545_9090 0.001
rdint_tsv2via_9_0 ndint_tsv_9_0 ndint_y_4545_909 0.001
rdint_tsv2via_9_2 ndint_tsv_9_2 ndint_y_4545_1818 0.001
rdint_tsv2via_9_4 ndint_tsv_9_4 ndint_y_4545_2727 0.001
rdint_tsv2via_9_6 ndint_tsv_9_6 ndint_y_4545_3636 0.001
rdint_tsv2via_9_8 ndint_tsv_9_8 ndint_y_4545_4545 0.001
rdint_tsv2via_9_10 ndint_tsv_9_10 ndint_xy_4545_5454 0.001
rdint_tsv2via_9_12 ndint_tsv_9_12 ndint_y_4545_6363 0.001
rdint_tsv2via_9_14 ndint_tsv_9_14 ndint_y_4545_7272 0.001
rdint_tsv2via_9_16 ndint_tsv_9_16 ndint_y_4545_8181 0.001
rdint_tsv2via_9_18 ndint_tsv_9_18 ndint_y_4545_9090 0.001
rdint_tsv2via_10_1 ndint_tsv_10_1 ndint_y_5454_909 0.001
rdint_tsv2via_10_3 ndint_tsv_10_3 ndint_y_5454_1818 0.001
rdint_tsv2via_10_5 ndint_tsv_10_5 ndint_y_5454_2727 0.001
rdint_tsv2via_10_7 ndint_tsv_10_7 ndint_y_5454_3636 0.001
rdint_tsv2via_10_9 ndint_tsv_10_9 ndint_xy_5454_4545 0.001
rdint_tsv2via_10_11 ndint_tsv_10_11 ndint_y_5454_5454 0.001
rdint_tsv2via_10_13 ndint_tsv_10_13 ndint_y_5454_6363 0.001
rdint_tsv2via_10_15 ndint_tsv_10_15 ndint_y_5454_7272 0.001
rdint_tsv2via_10_17 ndint_tsv_10_17 ndint_y_5454_8181 0.001
rdint_tsv2via_10_19 ndint_tsv_10_19 ndint_y_5454_9090 0.001
rdint_tsv2via_11_0 ndint_tsv_11_0 ndint_y_5454_909 0.001
rdint_tsv2via_11_2 ndint_tsv_11_2 ndint_y_5454_1818 0.001
rdint_tsv2via_11_4 ndint_tsv_11_4 ndint_y_5454_2727 0.001
rdint_tsv2via_11_6 ndint_tsv_11_6 ndint_y_5454_3636 0.001
rdint_tsv2via_11_8 ndint_tsv_11_8 ndint_xy_5454_4545 0.001
rdint_tsv2via_11_10 ndint_tsv_11_10 ndint_y_5454_5454 0.001
rdint_tsv2via_11_12 ndint_tsv_11_12 ndint_y_5454_6363 0.001
rdint_tsv2via_11_14 ndint_tsv_11_14 ndint_y_5454_7272 0.001
rdint_tsv2via_11_16 ndint_tsv_11_16 ndint_y_5454_8181 0.001
rdint_tsv2via_11_18 ndint_tsv_11_18 ndint_y_5454_9090 0.001
rdint_tsv2via_12_1 ndint_tsv_12_1 ndint_y_6363_909 0.001
rdint_tsv2via_12_3 ndint_tsv_12_3 ndint_y_6363_1818 0.001
rdint_tsv2via_12_5 ndint_tsv_12_5 ndint_y_6363_2727 0.001
rdint_tsv2via_12_7 ndint_tsv_12_7 ndint_xy_6363_3636 0.001
rdint_tsv2via_12_9 ndint_tsv_12_9 ndint_y_6363_4545 0.001
rdint_tsv2via_12_11 ndint_tsv_12_11 ndint_y_6363_5454 0.001
rdint_tsv2via_12_13 ndint_tsv_12_13 ndint_y_6363_6363 0.001
rdint_tsv2via_12_15 ndint_tsv_12_15 ndint_y_6363_7272 0.001
rdint_tsv2via_12_17 ndint_tsv_12_17 ndint_y_6363_8181 0.001
rdint_tsv2via_12_19 ndint_tsv_12_19 ndint_y_6363_9090 0.001
rdint_tsv2via_13_0 ndint_tsv_13_0 ndint_y_6363_909 0.001
rdint_tsv2via_13_2 ndint_tsv_13_2 ndint_y_6363_1818 0.001
rdint_tsv2via_13_4 ndint_tsv_13_4 ndint_y_6363_2727 0.001
rdint_tsv2via_13_6 ndint_tsv_13_6 ndint_xy_6363_3636 0.001
rdint_tsv2via_13_8 ndint_tsv_13_8 ndint_y_6363_4545 0.001
rdint_tsv2via_13_10 ndint_tsv_13_10 ndint_y_6363_5454 0.001
rdint_tsv2via_13_12 ndint_tsv_13_12 ndint_y_6363_6363 0.001
rdint_tsv2via_13_14 ndint_tsv_13_14 ndint_y_6363_7272 0.001
rdint_tsv2via_13_16 ndint_tsv_13_16 ndint_y_6363_8181 0.001
rdint_tsv2via_13_18 ndint_tsv_13_18 ndint_y_6363_9090 0.001
rdint_tsv2via_14_1 ndint_tsv_14_1 ndint_y_7272_909 0.001
rdint_tsv2via_14_3 ndint_tsv_14_3 ndint_y_7272_1818 0.001
rdint_tsv2via_14_5 ndint_tsv_14_5 ndint_xy_7272_2727 0.001
rdint_tsv2via_14_7 ndint_tsv_14_7 ndint_y_7272_3636 0.001
rdint_tsv2via_14_9 ndint_tsv_14_9 ndint_y_7272_4545 0.001
rdint_tsv2via_14_11 ndint_tsv_14_11 ndint_y_7272_5454 0.001
rdint_tsv2via_14_13 ndint_tsv_14_13 ndint_y_7272_6363 0.001
rdint_tsv2via_14_15 ndint_tsv_14_15 ndint_y_7272_7272 0.001
rdint_tsv2via_14_17 ndint_tsv_14_17 ndint_y_7272_8181 0.001
rdint_tsv2via_14_19 ndint_tsv_14_19 ndint_y_7272_9090 0.001
rdint_tsv2via_15_0 ndint_tsv_15_0 ndint_y_7272_909 0.001
rdint_tsv2via_15_2 ndint_tsv_15_2 ndint_y_7272_1818 0.001
rdint_tsv2via_15_4 ndint_tsv_15_4 ndint_xy_7272_2727 0.001
rdint_tsv2via_15_6 ndint_tsv_15_6 ndint_y_7272_3636 0.001
rdint_tsv2via_15_8 ndint_tsv_15_8 ndint_y_7272_4545 0.001
rdint_tsv2via_15_10 ndint_tsv_15_10 ndint_y_7272_5454 0.001
rdint_tsv2via_15_12 ndint_tsv_15_12 ndint_y_7272_6363 0.001
rdint_tsv2via_15_14 ndint_tsv_15_14 ndint_y_7272_7272 0.001
rdint_tsv2via_15_16 ndint_tsv_15_16 ndint_y_7272_8181 0.001
rdint_tsv2via_15_18 ndint_tsv_15_18 ndint_y_7272_9090 0.001
rdint_tsv2via_16_1 ndint_tsv_16_1 ndint_y_8181_909 0.001
rdint_tsv2via_16_3 ndint_tsv_16_3 ndint_xy_8181_1818 0.001
rdint_tsv2via_16_5 ndint_tsv_16_5 ndint_y_8181_2727 0.001
rdint_tsv2via_16_7 ndint_tsv_16_7 ndint_y_8181_3636 0.001
rdint_tsv2via_16_9 ndint_tsv_16_9 ndint_y_8181_4545 0.001
rdint_tsv2via_16_11 ndint_tsv_16_11 ndint_y_8181_5454 0.001
rdint_tsv2via_16_13 ndint_tsv_16_13 ndint_y_8181_6363 0.001
rdint_tsv2via_16_15 ndint_tsv_16_15 ndint_y_8181_7272 0.001
rdint_tsv2via_16_17 ndint_tsv_16_17 ndint_y_8181_8181 0.001
rdint_tsv2via_16_19 ndint_tsv_16_19 ndint_y_8181_9090 0.001
rdint_tsv2via_17_0 ndint_tsv_17_0 ndint_y_8181_909 0.001
rdint_tsv2via_17_2 ndint_tsv_17_2 ndint_xy_8181_1818 0.001
rdint_tsv2via_17_4 ndint_tsv_17_4 ndint_y_8181_2727 0.001
rdint_tsv2via_17_6 ndint_tsv_17_6 ndint_y_8181_3636 0.001
rdint_tsv2via_17_8 ndint_tsv_17_8 ndint_y_8181_4545 0.001
rdint_tsv2via_17_10 ndint_tsv_17_10 ndint_y_8181_5454 0.001
rdint_tsv2via_17_12 ndint_tsv_17_12 ndint_y_8181_6363 0.001
rdint_tsv2via_17_14 ndint_tsv_17_14 ndint_y_8181_7272 0.001
rdint_tsv2via_17_16 ndint_tsv_17_16 ndint_y_8181_8181 0.001
rdint_tsv2via_17_18 ndint_tsv_17_18 ndint_y_8181_9090 0.001
rdint_tsv2via_18_1 ndint_tsv_18_1 ndint_xy_9090_909 0.001
rdint_tsv2via_18_3 ndint_tsv_18_3 ndint_y_9090_1818 0.001
rdint_tsv2via_18_5 ndint_tsv_18_5 ndint_y_9090_2727 0.001
rdint_tsv2via_18_7 ndint_tsv_18_7 ndint_y_9090_3636 0.001
rdint_tsv2via_18_9 ndint_tsv_18_9 ndint_y_9090_4545 0.001
rdint_tsv2via_18_11 ndint_tsv_18_11 ndint_y_9090_5454 0.001
rdint_tsv2via_18_13 ndint_tsv_18_13 ndint_y_9090_6363 0.001
rdint_tsv2via_18_15 ndint_tsv_18_15 ndint_y_9090_7272 0.001
rdint_tsv2via_18_17 ndint_tsv_18_17 ndint_y_9090_8181 0.001
rdint_tsv2via_18_19 ndint_tsv_18_19 ndint_y_9090_9090 0.001
rdint_tsv2via_19_0 ndint_tsv_19_0 ndint_xy_9090_909 0.001
rdint_tsv2via_19_2 ndint_tsv_19_2 ndint_y_9090_1818 0.001
rdint_tsv2via_19_4 ndint_tsv_19_4 ndint_y_9090_2727 0.001
rdint_tsv2via_19_6 ndint_tsv_19_6 ndint_y_9090_3636 0.001
rdint_tsv2via_19_8 ndint_tsv_19_8 ndint_y_9090_4545 0.001
rdint_tsv2via_19_10 ndint_tsv_19_10 ndint_y_9090_5454 0.001
rdint_tsv2via_19_12 ndint_tsv_19_12 ndint_y_9090_6363 0.001
rdint_tsv2via_19_14 ndint_tsv_19_14 ndint_y_9090_7272 0.001
rdint_tsv2via_19_16 ndint_tsv_19_16 ndint_y_9090_8181 0.001
rdint_tsv2via_19_18 ndint_tsv_19_18 ndint_y_9090_9090 0.001

*-- tsv bump array to pkg
rdint_tsv_0_1 ndint_bump_0_1 nd_pkg_pad 0.001
rdint_tsv_0_3 ndint_bump_0_3 nd_pkg_pad 0.001
rdint_tsv_0_5 ndint_bump_0_5 nd_pkg_pad 0.001
rdint_tsv_0_7 ndint_bump_0_7 nd_pkg_pad 0.001
rdint_tsv_0_9 ndint_bump_0_9 nd_pkg_pad 0.001
rdint_tsv_0_11 ndint_bump_0_11 nd_pkg_pad 0.001
rdint_tsv_0_13 ndint_bump_0_13 nd_pkg_pad 0.001
rdint_tsv_0_15 ndint_bump_0_15 nd_pkg_pad 0.001
rdint_tsv_0_17 ndint_bump_0_17 nd_pkg_pad 0.001
rdint_tsv_0_19 ndint_bump_0_19 nd_pkg_pad 0.001
rdint_tsv_1_0 ndint_bump_1_0 nd_pkg_pad 0.001
rdint_tsv_1_2 ndint_bump_1_2 nd_pkg_pad 0.001
rdint_tsv_1_4 ndint_bump_1_4 nd_pkg_pad 0.001
rdint_tsv_1_6 ndint_bump_1_6 nd_pkg_pad 0.001
rdint_tsv_1_8 ndint_bump_1_8 nd_pkg_pad 0.001
rdint_tsv_1_10 ndint_bump_1_10 nd_pkg_pad 0.001
rdint_tsv_1_12 ndint_bump_1_12 nd_pkg_pad 0.001
rdint_tsv_1_14 ndint_bump_1_14 nd_pkg_pad 0.001
rdint_tsv_1_16 ndint_bump_1_16 nd_pkg_pad 0.001
rdint_tsv_1_18 ndint_bump_1_18 nd_pkg_pad 0.001
rdint_tsv_2_1 ndint_bump_2_1 nd_pkg_pad 0.001
rdint_tsv_2_3 ndint_bump_2_3 nd_pkg_pad 0.001
rdint_tsv_2_5 ndint_bump_2_5 nd_pkg_pad 0.001
rdint_tsv_2_7 ndint_bump_2_7 nd_pkg_pad 0.001
rdint_tsv_2_9 ndint_bump_2_9 nd_pkg_pad 0.001
rdint_tsv_2_11 ndint_bump_2_11 nd_pkg_pad 0.001
rdint_tsv_2_13 ndint_bump_2_13 nd_pkg_pad 0.001
rdint_tsv_2_15 ndint_bump_2_15 nd_pkg_pad 0.001
rdint_tsv_2_17 ndint_bump_2_17 nd_pkg_pad 0.001
rdint_tsv_2_19 ndint_bump_2_19 nd_pkg_pad 0.001
rdint_tsv_3_0 ndint_bump_3_0 nd_pkg_pad 0.001
rdint_tsv_3_2 ndint_bump_3_2 nd_pkg_pad 0.001
rdint_tsv_3_4 ndint_bump_3_4 nd_pkg_pad 0.001
rdint_tsv_3_6 ndint_bump_3_6 nd_pkg_pad 0.001
rdint_tsv_3_8 ndint_bump_3_8 nd_pkg_pad 0.001
rdint_tsv_3_10 ndint_bump_3_10 nd_pkg_pad 0.001
rdint_tsv_3_12 ndint_bump_3_12 nd_pkg_pad 0.001
rdint_tsv_3_14 ndint_bump_3_14 nd_pkg_pad 0.001
rdint_tsv_3_16 ndint_bump_3_16 nd_pkg_pad 0.001
rdint_tsv_3_18 ndint_bump_3_18 nd_pkg_pad 0.001
rdint_tsv_4_1 ndint_bump_4_1 nd_pkg_pad 0.001
rdint_tsv_4_3 ndint_bump_4_3 nd_pkg_pad 0.001
rdint_tsv_4_5 ndint_bump_4_5 nd_pkg_pad 0.001
rdint_tsv_4_7 ndint_bump_4_7 nd_pkg_pad 0.001
rdint_tsv_4_9 ndint_bump_4_9 nd_pkg_pad 0.001
rdint_tsv_4_11 ndint_bump_4_11 nd_pkg_pad 0.001
rdint_tsv_4_13 ndint_bump_4_13 nd_pkg_pad 0.001
rdint_tsv_4_15 ndint_bump_4_15 nd_pkg_pad 0.001
rdint_tsv_4_17 ndint_bump_4_17 nd_pkg_pad 0.001
rdint_tsv_4_19 ndint_bump_4_19 nd_pkg_pad 0.001
rdint_tsv_5_0 ndint_bump_5_0 nd_pkg_pad 0.001
rdint_tsv_5_2 ndint_bump_5_2 nd_pkg_pad 0.001
rdint_tsv_5_4 ndint_bump_5_4 nd_pkg_pad 0.001
rdint_tsv_5_6 ndint_bump_5_6 nd_pkg_pad 0.001
rdint_tsv_5_8 ndint_bump_5_8 nd_pkg_pad 0.001
rdint_tsv_5_10 ndint_bump_5_10 nd_pkg_pad 0.001
rdint_tsv_5_12 ndint_bump_5_12 nd_pkg_pad 0.001
rdint_tsv_5_14 ndint_bump_5_14 nd_pkg_pad 0.001
rdint_tsv_5_16 ndint_bump_5_16 nd_pkg_pad 0.001
rdint_tsv_5_18 ndint_bump_5_18 nd_pkg_pad 0.001
rdint_tsv_6_1 ndint_bump_6_1 nd_pkg_pad 0.001
rdint_tsv_6_3 ndint_bump_6_3 nd_pkg_pad 0.001
rdint_tsv_6_5 ndint_bump_6_5 nd_pkg_pad 0.001
rdint_tsv_6_7 ndint_bump_6_7 nd_pkg_pad 0.001
rdint_tsv_6_9 ndint_bump_6_9 nd_pkg_pad 0.001
rdint_tsv_6_11 ndint_bump_6_11 nd_pkg_pad 0.001
rdint_tsv_6_13 ndint_bump_6_13 nd_pkg_pad 0.001
rdint_tsv_6_15 ndint_bump_6_15 nd_pkg_pad 0.001
rdint_tsv_6_17 ndint_bump_6_17 nd_pkg_pad 0.001
rdint_tsv_6_19 ndint_bump_6_19 nd_pkg_pad 0.001
rdint_tsv_7_0 ndint_bump_7_0 nd_pkg_pad 0.001
rdint_tsv_7_2 ndint_bump_7_2 nd_pkg_pad 0.001
rdint_tsv_7_4 ndint_bump_7_4 nd_pkg_pad 0.001
rdint_tsv_7_6 ndint_bump_7_6 nd_pkg_pad 0.001
rdint_tsv_7_8 ndint_bump_7_8 nd_pkg_pad 0.001
rdint_tsv_7_10 ndint_bump_7_10 nd_pkg_pad 0.001
rdint_tsv_7_12 ndint_bump_7_12 nd_pkg_pad 0.001
rdint_tsv_7_14 ndint_bump_7_14 nd_pkg_pad 0.001
rdint_tsv_7_16 ndint_bump_7_16 nd_pkg_pad 0.001
rdint_tsv_7_18 ndint_bump_7_18 nd_pkg_pad 0.001
rdint_tsv_8_1 ndint_bump_8_1 nd_pkg_pad 0.001
rdint_tsv_8_3 ndint_bump_8_3 nd_pkg_pad 0.001
rdint_tsv_8_5 ndint_bump_8_5 nd_pkg_pad 0.001
rdint_tsv_8_7 ndint_bump_8_7 nd_pkg_pad 0.001
rdint_tsv_8_9 ndint_bump_8_9 nd_pkg_pad 0.001
rdint_tsv_8_11 ndint_bump_8_11 nd_pkg_pad 0.001
rdint_tsv_8_13 ndint_bump_8_13 nd_pkg_pad 0.001
rdint_tsv_8_15 ndint_bump_8_15 nd_pkg_pad 0.001
rdint_tsv_8_17 ndint_bump_8_17 nd_pkg_pad 0.001
rdint_tsv_8_19 ndint_bump_8_19 nd_pkg_pad 0.001
rdint_tsv_9_0 ndint_bump_9_0 nd_pkg_pad 0.001
rdint_tsv_9_2 ndint_bump_9_2 nd_pkg_pad 0.001
rdint_tsv_9_4 ndint_bump_9_4 nd_pkg_pad 0.001
rdint_tsv_9_6 ndint_bump_9_6 nd_pkg_pad 0.001
rdint_tsv_9_8 ndint_bump_9_8 nd_pkg_pad 0.001
rdint_tsv_9_10 ndint_bump_9_10 nd_pkg_pad 0.001
rdint_tsv_9_12 ndint_bump_9_12 nd_pkg_pad 0.001
rdint_tsv_9_14 ndint_bump_9_14 nd_pkg_pad 0.001
rdint_tsv_9_16 ndint_bump_9_16 nd_pkg_pad 0.001
rdint_tsv_9_18 ndint_bump_9_18 nd_pkg_pad 0.001
rdint_tsv_10_1 ndint_bump_10_1 nd_pkg_pad 0.001
rdint_tsv_10_3 ndint_bump_10_3 nd_pkg_pad 0.001
rdint_tsv_10_5 ndint_bump_10_5 nd_pkg_pad 0.001
rdint_tsv_10_7 ndint_bump_10_7 nd_pkg_pad 0.001
rdint_tsv_10_9 ndint_bump_10_9 nd_pkg_pad 0.001
rdint_tsv_10_11 ndint_bump_10_11 nd_pkg_pad 0.001
rdint_tsv_10_13 ndint_bump_10_13 nd_pkg_pad 0.001
rdint_tsv_10_15 ndint_bump_10_15 nd_pkg_pad 0.001
rdint_tsv_10_17 ndint_bump_10_17 nd_pkg_pad 0.001
rdint_tsv_10_19 ndint_bump_10_19 nd_pkg_pad 0.001
rdint_tsv_11_0 ndint_bump_11_0 nd_pkg_pad 0.001
rdint_tsv_11_2 ndint_bump_11_2 nd_pkg_pad 0.001
rdint_tsv_11_4 ndint_bump_11_4 nd_pkg_pad 0.001
rdint_tsv_11_6 ndint_bump_11_6 nd_pkg_pad 0.001
rdint_tsv_11_8 ndint_bump_11_8 nd_pkg_pad 0.001
rdint_tsv_11_10 ndint_bump_11_10 nd_pkg_pad 0.001
rdint_tsv_11_12 ndint_bump_11_12 nd_pkg_pad 0.001
rdint_tsv_11_14 ndint_bump_11_14 nd_pkg_pad 0.001
rdint_tsv_11_16 ndint_bump_11_16 nd_pkg_pad 0.001
rdint_tsv_11_18 ndint_bump_11_18 nd_pkg_pad 0.001
rdint_tsv_12_1 ndint_bump_12_1 nd_pkg_pad 0.001
rdint_tsv_12_3 ndint_bump_12_3 nd_pkg_pad 0.001
rdint_tsv_12_5 ndint_bump_12_5 nd_pkg_pad 0.001
rdint_tsv_12_7 ndint_bump_12_7 nd_pkg_pad 0.001
rdint_tsv_12_9 ndint_bump_12_9 nd_pkg_pad 0.001
rdint_tsv_12_11 ndint_bump_12_11 nd_pkg_pad 0.001
rdint_tsv_12_13 ndint_bump_12_13 nd_pkg_pad 0.001
rdint_tsv_12_15 ndint_bump_12_15 nd_pkg_pad 0.001
rdint_tsv_12_17 ndint_bump_12_17 nd_pkg_pad 0.001
rdint_tsv_12_19 ndint_bump_12_19 nd_pkg_pad 0.001
rdint_tsv_13_0 ndint_bump_13_0 nd_pkg_pad 0.001
rdint_tsv_13_2 ndint_bump_13_2 nd_pkg_pad 0.001
rdint_tsv_13_4 ndint_bump_13_4 nd_pkg_pad 0.001
rdint_tsv_13_6 ndint_bump_13_6 nd_pkg_pad 0.001
rdint_tsv_13_8 ndint_bump_13_8 nd_pkg_pad 0.001
rdint_tsv_13_10 ndint_bump_13_10 nd_pkg_pad 0.001
rdint_tsv_13_12 ndint_bump_13_12 nd_pkg_pad 0.001
rdint_tsv_13_14 ndint_bump_13_14 nd_pkg_pad 0.001
rdint_tsv_13_16 ndint_bump_13_16 nd_pkg_pad 0.001
rdint_tsv_13_18 ndint_bump_13_18 nd_pkg_pad 0.001
rdint_tsv_14_1 ndint_bump_14_1 nd_pkg_pad 0.001
rdint_tsv_14_3 ndint_bump_14_3 nd_pkg_pad 0.001
rdint_tsv_14_5 ndint_bump_14_5 nd_pkg_pad 0.001
rdint_tsv_14_7 ndint_bump_14_7 nd_pkg_pad 0.001
rdint_tsv_14_9 ndint_bump_14_9 nd_pkg_pad 0.001
rdint_tsv_14_11 ndint_bump_14_11 nd_pkg_pad 0.001
rdint_tsv_14_13 ndint_bump_14_13 nd_pkg_pad 0.001
rdint_tsv_14_15 ndint_bump_14_15 nd_pkg_pad 0.001
rdint_tsv_14_17 ndint_bump_14_17 nd_pkg_pad 0.001
rdint_tsv_14_19 ndint_bump_14_19 nd_pkg_pad 0.001
rdint_tsv_15_0 ndint_bump_15_0 nd_pkg_pad 0.001
rdint_tsv_15_2 ndint_bump_15_2 nd_pkg_pad 0.001
rdint_tsv_15_4 ndint_bump_15_4 nd_pkg_pad 0.001
rdint_tsv_15_6 ndint_bump_15_6 nd_pkg_pad 0.001
rdint_tsv_15_8 ndint_bump_15_8 nd_pkg_pad 0.001
rdint_tsv_15_10 ndint_bump_15_10 nd_pkg_pad 0.001
rdint_tsv_15_12 ndint_bump_15_12 nd_pkg_pad 0.001
rdint_tsv_15_14 ndint_bump_15_14 nd_pkg_pad 0.001
rdint_tsv_15_16 ndint_bump_15_16 nd_pkg_pad 0.001
rdint_tsv_15_18 ndint_bump_15_18 nd_pkg_pad 0.001
rdint_tsv_16_1 ndint_bump_16_1 nd_pkg_pad 0.001
rdint_tsv_16_3 ndint_bump_16_3 nd_pkg_pad 0.001
rdint_tsv_16_5 ndint_bump_16_5 nd_pkg_pad 0.001
rdint_tsv_16_7 ndint_bump_16_7 nd_pkg_pad 0.001
rdint_tsv_16_9 ndint_bump_16_9 nd_pkg_pad 0.001
rdint_tsv_16_11 ndint_bump_16_11 nd_pkg_pad 0.001
rdint_tsv_16_13 ndint_bump_16_13 nd_pkg_pad 0.001
rdint_tsv_16_15 ndint_bump_16_15 nd_pkg_pad 0.001
rdint_tsv_16_17 ndint_bump_16_17 nd_pkg_pad 0.001
rdint_tsv_16_19 ndint_bump_16_19 nd_pkg_pad 0.001
rdint_tsv_17_0 ndint_bump_17_0 nd_pkg_pad 0.001
rdint_tsv_17_2 ndint_bump_17_2 nd_pkg_pad 0.001
rdint_tsv_17_4 ndint_bump_17_4 nd_pkg_pad 0.001
rdint_tsv_17_6 ndint_bump_17_6 nd_pkg_pad 0.001
rdint_tsv_17_8 ndint_bump_17_8 nd_pkg_pad 0.001
rdint_tsv_17_10 ndint_bump_17_10 nd_pkg_pad 0.001
rdint_tsv_17_12 ndint_bump_17_12 nd_pkg_pad 0.001
rdint_tsv_17_14 ndint_bump_17_14 nd_pkg_pad 0.001
rdint_tsv_17_16 ndint_bump_17_16 nd_pkg_pad 0.001
rdint_tsv_17_18 ndint_bump_17_18 nd_pkg_pad 0.001
rdint_tsv_18_1 ndint_bump_18_1 nd_pkg_pad 0.001
rdint_tsv_18_3 ndint_bump_18_3 nd_pkg_pad 0.001
rdint_tsv_18_5 ndint_bump_18_5 nd_pkg_pad 0.001
rdint_tsv_18_7 ndint_bump_18_7 nd_pkg_pad 0.001
rdint_tsv_18_9 ndint_bump_18_9 nd_pkg_pad 0.001
rdint_tsv_18_11 ndint_bump_18_11 nd_pkg_pad 0.001
rdint_tsv_18_13 ndint_bump_18_13 nd_pkg_pad 0.001
rdint_tsv_18_15 ndint_bump_18_15 nd_pkg_pad 0.001
rdint_tsv_18_17 ndint_bump_18_17 nd_pkg_pad 0.001
rdint_tsv_18_19 ndint_bump_18_19 nd_pkg_pad 0.001
rdint_tsv_19_0 ndint_bump_19_0 nd_pkg_pad 0.001
rdint_tsv_19_2 ndint_bump_19_2 nd_pkg_pad 0.001
rdint_tsv_19_4 ndint_bump_19_4 nd_pkg_pad 0.001
rdint_tsv_19_6 ndint_bump_19_6 nd_pkg_pad 0.001
rdint_tsv_19_8 ndint_bump_19_8 nd_pkg_pad 0.001
rdint_tsv_19_10 ndint_bump_19_10 nd_pkg_pad 0.001
rdint_tsv_19_12 ndint_bump_19_12 nd_pkg_pad 0.001
rdint_tsv_19_14 ndint_bump_19_14 nd_pkg_pad 0.001
rdint_tsv_19_16 ndint_bump_19_16 nd_pkg_pad 0.001
rdint_tsv_19_18 ndint_bump_19_18 nd_pkg_pad 0.001

*-- pkg instances
xpkg_vdd vdd_pkg nd_pkg_pad pkg_model
xpkg_vss vss_pkg ns_pkg_pad pkg_model
.include 'pkg.subckt'

*-- pcb instances
xpcb_vdd vdd vdd_pkg pcb_model
xpcb_vss vss vss_pkg pcb_model
.include 'pcb.subckt'


*-- external power source
ivdd 0 vdd 0 ac 1
ivss 0 vss 0 ac 1
.ac dec 100 1e+06 1e+10
.end
